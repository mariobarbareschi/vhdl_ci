----------------------------------------------------------------------------------
-- Engineer: 		Marcello Traiola
--
-- Create Date: 9:59:52 20/10/2017
-- Design Name: 
-- Module Name: 
-- Project Name: 
-- Revision 1.0 - File Created
-- Notes - File generated using XbarGen tool by Marcello Traiola (marcellotraiola@gmail.com)
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library memristor_lib;
use memristor_lib.types.all;

use work.crossbar_structure_1.all;

entity crossbar_controller_1 is
Port ( 
pi26 : in  STD_LOGIC;
pi15 : in  STD_LOGIC;
lo6 : in  STD_LOGIC;
lo5 : in  STD_LOGIC;
lo4 : in  STD_LOGIC;
lo3 : in  STD_LOGIC;
lo2 : in  STD_LOGIC;
lo1 : in  STD_LOGIC;
lo0 : in  STD_LOGIC;
pi00 : in  STD_LOGIC;
pi06 : in  STD_LOGIC;
pi03 : in  STD_LOGIC;
pi07 : in  STD_LOGIC;
pi08 : in  STD_LOGIC;
pi09 : in  STD_LOGIC;
pi10 : in  STD_LOGIC;
pi02 : in  STD_LOGIC;
pi17 : in  STD_LOGIC;
pi01 : in  STD_LOGIC;
pi11 : in  STD_LOGIC;
pi12 : in  STD_LOGIC;
pi13 : in  STD_LOGIC;
pi14 : in  STD_LOGIC;
pi04 : in  STD_LOGIC;
pi16 : in  STD_LOGIC;
pi05 : in  STD_LOGIC;
pi18 : in  STD_LOGIC;
pi19 : in  STD_LOGIC;
pi20 : in  STD_LOGIC;
pi21 : in  STD_LOGIC;
pi22 : in  STD_LOGIC;
pi23 : in  STD_LOGIC;
pi24 : in  STD_LOGIC;
pi25 : in  STD_LOGIC;
en : in STD_LOGIC;
po00 : out  STD_LOGIC;
po01 : out  STD_LOGIC;
po02 : out  STD_LOGIC;
po03 : out  STD_LOGIC;
po04 : out  STD_LOGIC;
po05 : out  STD_LOGIC;
po06 : out  STD_LOGIC;
po07 : out  STD_LOGIC;
po08 : out  STD_LOGIC;
po09 : out  STD_LOGIC;
po10 : out  STD_LOGIC;
po11 : out  STD_LOGIC;
po12 : out  STD_LOGIC;
po13 : out  STD_LOGIC;
po15 : out  STD_LOGIC;
po16 : out  STD_LOGIC;
po17 : out  STD_LOGIC;
po18 : out  STD_LOGIC;
po20 : out  STD_LOGIC;
po21 : out  STD_LOGIC;
po22 : out  STD_LOGIC;
po23 : out  STD_LOGIC;
po24 : out  STD_LOGIC;
po25 : out  STD_LOGIC;
po26 : out  STD_LOGIC;
po27 : out  STD_LOGIC;
po28 : out  STD_LOGIC;
po29 : out  STD_LOGIC;
po30 : out  STD_LOGIC;
po31 : out  STD_LOGIC;
po32 : out  STD_LOGIC;
po33 : out  STD_LOGIC;
po34 : out  STD_LOGIC;
po35 : out  STD_LOGIC;
po36 : out  STD_LOGIC;
po37 : out  STD_LOGIC;
po38 : out  STD_LOGIC;
po39 : out  STD_LOGIC;
po40 : out  STD_LOGIC;
po41 : out  STD_LOGIC;
po42 : out  STD_LOGIC;
po43 : out  STD_LOGIC;
po44 : out  STD_LOGIC;
po45 : out  STD_LOGIC;
po46 : out  STD_LOGIC;
po47 : out  STD_LOGIC;
po48 : out  STD_LOGIC;
po49 : out  STD_LOGIC;
po50 : out  STD_LOGIC;
po51 : out  STD_LOGIC;
po52 : out  STD_LOGIC;
po53 : out  STD_LOGIC;
po54 : out  STD_LOGIC;
po55 : out  STD_LOGIC;
li0 : out  STD_LOGIC;
li1 : out  STD_LOGIC;
li2 : out  STD_LOGIC;
li3 : out  STD_LOGIC;
li4 : out  STD_LOGIC;
li5 : out  STD_LOGIC;
li6 : out  STD_LOGIC;
done : out STD_LOGIC
);
end crossbar_controller_1;

architecture Behavioral of crossbar_controller_1 is

COMPONENT crossbar_1
PORT(
Vpos : IN voltage_vector(0 to 189);
Vneg : IN voltage_vector(0 to 735);
output : out STD_LOGIC_VECTOR(0 to 60) --here we have 61 outputs
);
END COMPONENT;

signal Vpos_temp : voltage_vector(0 to 189);
signal Vneg_temp: voltage_vector(0 to 735);
signal output_temp : STD_LOGIC_VECTOR(0 to 60);

	alias XbG_V0 : voltage is Vpos_temp(0);
	alias XbG_V1 : voltage is Vpos_temp(1);
	alias XbG_V2 : voltage is Vpos_temp(2);
	alias XbG_V3 : voltage is Vpos_temp(3);
	alias XbG_V4 : voltage is Vpos_temp(4);
	alias XbG_V5 : voltage is Vpos_temp(5);
	alias XbG_V6 : voltage is Vpos_temp(6);
	alias XbG_V7 : voltage is Vpos_temp(7);
	alias XbG_V8 : voltage is Vpos_temp(8);
	alias XbG_V9 : voltage is Vpos_temp(9);
	alias XbG_V10 : voltage is Vpos_temp(10);
	alias XbG_V11 : voltage is Vpos_temp(11);
	alias XbG_V12 : voltage is Vpos_temp(12);
	alias XbG_V13 : voltage is Vpos_temp(13);
	alias XbG_V14 : voltage is Vpos_temp(14);
	alias XbG_V15 : voltage is Vpos_temp(15);
	alias XbG_V16 : voltage is Vpos_temp(16);
	alias XbG_V17 : voltage is Vpos_temp(17);
	alias XbG_V18 : voltage is Vpos_temp(18);
	alias XbG_V19 : voltage is Vpos_temp(19);
	alias XbG_V20 : voltage is Vpos_temp(20);
	alias XbG_V21 : voltage is Vpos_temp(21);
	alias XbG_V22 : voltage is Vpos_temp(22);
	alias XbG_V23 : voltage is Vpos_temp(23);
	alias XbG_V24 : voltage is Vpos_temp(24);
	alias XbG_V25 : voltage is Vpos_temp(25);
	alias XbG_V26 : voltage is Vpos_temp(26);
	alias XbG_V27 : voltage is Vpos_temp(27);
	alias XbG_V28 : voltage is Vpos_temp(28);
	alias XbG_V29 : voltage is Vpos_temp(29);
	alias XbG_V30 : voltage is Vpos_temp(30);
	alias XbG_V31 : voltage is Vpos_temp(31);
	alias XbG_V32 : voltage is Vpos_temp(32);
	alias XbG_V33 : voltage is Vpos_temp(33);
	alias XbG_V34 : voltage is Vpos_temp(34);
	alias XbG_V35 : voltage is Vpos_temp(35);
	alias XbG_V36 : voltage is Vpos_temp(36);
	alias XbG_V37 : voltage is Vpos_temp(37);
	alias XbG_V38 : voltage is Vpos_temp(38);
	alias XbG_V39 : voltage is Vpos_temp(39);
	alias XbG_V40 : voltage is Vpos_temp(40);
	alias XbG_V41 : voltage is Vpos_temp(41);
	alias XbG_V42 : voltage is Vpos_temp(42);
	alias XbG_V43 : voltage is Vpos_temp(43);
	alias XbG_V44 : voltage is Vpos_temp(44);
	alias XbG_V45 : voltage is Vpos_temp(45);
	alias XbG_V46 : voltage is Vpos_temp(46);
	alias XbG_V47 : voltage is Vpos_temp(47);
	alias XbG_V48 : voltage is Vpos_temp(48);
	alias XbG_V49 : voltage is Vpos_temp(49);
	alias XbG_V50 : voltage is Vpos_temp(50);
	alias XbG_V51 : voltage is Vpos_temp(51);
	alias XbG_V52 : voltage is Vpos_temp(52);
	alias XbG_V53 : voltage is Vpos_temp(53);
	alias XbG_V54 : voltage is Vpos_temp(54);
	alias XbG_V55 : voltage is Vpos_temp(55);
	alias XbG_V56 : voltage is Vpos_temp(56);
	alias XbG_V57 : voltage is Vpos_temp(57);
	alias XbG_V58 : voltage is Vpos_temp(58);
	alias XbG_V59 : voltage is Vpos_temp(59);
	alias XbG_V60 : voltage is Vpos_temp(60);
	alias XbG_V61 : voltage is Vpos_temp(61);
	alias XbG_V62 : voltage is Vpos_temp(62);
	alias XbG_V63 : voltage is Vpos_temp(63);
	alias XbG_V64 : voltage is Vpos_temp(64);
	alias XbG_V65 : voltage is Vpos_temp(65);
	alias XbG_V66 : voltage is Vpos_temp(66);
	alias XbG_V67 : voltage is Vpos_temp(67);
	alias XbG_V68 : voltage is Vpos_temp(68);
	alias XbG_V69 : voltage is Vpos_temp(69);
	alias XbG_V70 : voltage is Vpos_temp(70);
	alias XbG_V71 : voltage is Vpos_temp(71);
	alias XbG_V72 : voltage is Vpos_temp(72);
	alias XbG_V73 : voltage is Vpos_temp(73);
	alias XbG_V74 : voltage is Vpos_temp(74);
	alias XbG_V75 : voltage is Vpos_temp(75);
	alias XbG_V76 : voltage is Vpos_temp(76);
	alias XbG_V77 : voltage is Vpos_temp(77);
	alias XbG_V78 : voltage is Vpos_temp(78);
	alias XbG_V79 : voltage is Vpos_temp(79);
	alias XbG_V80 : voltage is Vpos_temp(80);
	alias XbG_V81 : voltage is Vpos_temp(81);
	alias XbG_V82 : voltage is Vpos_temp(82);
	alias XbG_V83 : voltage is Vpos_temp(83);
	alias XbG_V84 : voltage is Vpos_temp(84);
	alias XbG_V85 : voltage is Vpos_temp(85);
	alias XbG_V86 : voltage is Vpos_temp(86);
	alias XbG_V87 : voltage is Vpos_temp(87);
	alias XbG_V88 : voltage is Vpos_temp(88);
	alias XbG_V89 : voltage is Vpos_temp(89);
	alias XbG_V90 : voltage is Vpos_temp(90);
	alias XbG_V91 : voltage is Vpos_temp(91);
	alias XbG_V92 : voltage is Vpos_temp(92);
	alias XbG_V93 : voltage is Vpos_temp(93);
	alias XbG_V94 : voltage is Vpos_temp(94);
	alias XbG_V95 : voltage is Vpos_temp(95);
	alias XbG_V96 : voltage is Vpos_temp(96);
	alias XbG_V97 : voltage is Vpos_temp(97);
	alias XbG_V98 : voltage is Vpos_temp(98);
	alias XbG_V99 : voltage is Vpos_temp(99);
	alias XbG_V100 : voltage is Vpos_temp(100);
	alias XbG_V101 : voltage is Vpos_temp(101);
	alias XbG_V102 : voltage is Vpos_temp(102);
	alias XbG_V103 : voltage is Vpos_temp(103);
	alias XbG_V104 : voltage is Vpos_temp(104);
	alias XbG_V105 : voltage is Vpos_temp(105);
	alias XbG_V106 : voltage is Vpos_temp(106);
	alias XbG_V107 : voltage is Vpos_temp(107);
	alias XbG_V108 : voltage is Vpos_temp(108);
	alias XbG_V109 : voltage is Vpos_temp(109);
	alias XbG_V110 : voltage is Vpos_temp(110);
	alias XbG_V111 : voltage is Vpos_temp(111);
	alias XbG_V112 : voltage is Vpos_temp(112);
	alias XbG_V113 : voltage is Vpos_temp(113);
	alias XbG_V114 : voltage is Vpos_temp(114);
	alias XbG_V115 : voltage is Vpos_temp(115);
	alias XbG_V116 : voltage is Vpos_temp(116);
	alias XbG_V117 : voltage is Vpos_temp(117);
	alias XbG_V118 : voltage is Vpos_temp(118);
	alias XbG_V119 : voltage is Vpos_temp(119);
	alias XbG_V120 : voltage is Vpos_temp(120);
	alias XbG_V121 : voltage is Vpos_temp(121);
	alias XbG_V122 : voltage is Vpos_temp(122);
	alias XbG_V123 : voltage is Vpos_temp(123);
	alias XbG_V124 : voltage is Vpos_temp(124);
	alias XbG_V125 : voltage is Vpos_temp(125);
	alias XbG_V126 : voltage is Vpos_temp(126);
	alias XbG_V127 : voltage is Vpos_temp(127);
	alias XbG_V128 : voltage is Vpos_temp(128);
	alias XbG_V129 : voltage is Vpos_temp(129);
	alias XbG_V130 : voltage is Vpos_temp(130);
	alias XbG_V131 : voltage is Vpos_temp(131);
	alias XbG_V132 : voltage is Vpos_temp(132);
	alias XbG_V133 : voltage is Vpos_temp(133);
	alias XbG_V134 : voltage is Vpos_temp(134);
	alias XbG_V135 : voltage is Vpos_temp(135);
	alias XbG_V136 : voltage is Vpos_temp(136);
	alias XbG_V137 : voltage is Vpos_temp(137);
	alias XbG_V138 : voltage is Vpos_temp(138);
	alias XbG_V139 : voltage is Vpos_temp(139);
	alias XbG_V140 : voltage is Vpos_temp(140);
	alias XbG_V141 : voltage is Vpos_temp(141);
	alias XbG_V142 : voltage is Vpos_temp(142);
	alias XbG_V143 : voltage is Vpos_temp(143);
	alias XbG_V144 : voltage is Vpos_temp(144);
	alias XbG_V145 : voltage is Vpos_temp(145);
	alias XbG_V146 : voltage is Vpos_temp(146);
	alias XbG_V147 : voltage is Vpos_temp(147);
	alias XbG_V148 : voltage is Vpos_temp(148);
	alias XbG_V149 : voltage is Vpos_temp(149);
	alias XbG_V150 : voltage is Vpos_temp(150);
	alias XbG_V151 : voltage is Vpos_temp(151);
	alias XbG_V152 : voltage is Vpos_temp(152);
	alias XbG_V153 : voltage is Vpos_temp(153);
	alias XbG_V154 : voltage is Vpos_temp(154);
	alias XbG_V155 : voltage is Vpos_temp(155);
	alias XbG_V156 : voltage is Vpos_temp(156);
	alias XbG_V157 : voltage is Vpos_temp(157);
	alias XbG_V158 : voltage is Vpos_temp(158);
	alias XbG_V159 : voltage is Vpos_temp(159);
	alias XbG_V160 : voltage is Vpos_temp(160);
	alias XbG_V161 : voltage is Vpos_temp(161);
	alias XbG_V162 : voltage is Vpos_temp(162);
	alias XbG_V163 : voltage is Vpos_temp(163);
	alias XbG_V164 : voltage is Vpos_temp(164);
	alias XbG_V165 : voltage is Vpos_temp(165);
	alias XbG_V166 : voltage is Vpos_temp(166);
	alias XbG_V167 : voltage is Vpos_temp(167);
	alias XbG_V168 : voltage is Vpos_temp(168);
	alias XbG_V169 : voltage is Vpos_temp(169);
	alias XbG_V170 : voltage is Vpos_temp(170);
	alias XbG_V171 : voltage is Vpos_temp(171);
	alias XbG_V172 : voltage is Vpos_temp(172);
	alias XbG_V173 : voltage is Vpos_temp(173);
	alias XbG_V174 : voltage is Vpos_temp(174);
	alias XbG_V175 : voltage is Vpos_temp(175);
	alias XbG_V176 : voltage is Vpos_temp(176);
	alias XbG_V177 : voltage is Vpos_temp(177);
	alias XbG_V178 : voltage is Vpos_temp(178);
	alias XbG_V179 : voltage is Vpos_temp(179);
	alias XbG_V180 : voltage is Vpos_temp(180);
	alias XbG_V181 : voltage is Vpos_temp(181);
	alias XbG_V182 : voltage is Vpos_temp(182);
	alias XbG_V183 : voltage is Vpos_temp(183);
	alias XbG_V184 : voltage is Vpos_temp(184);
	alias XbG_V185 : voltage is Vpos_temp(185);
	alias XbG_V186 : voltage is Vpos_temp(186);
	alias XbG_V187 : voltage is Vpos_temp(187);
	alias XbG_V188 : voltage is Vpos_temp(188);
	alias XbG_V189 : voltage is Vpos_temp(189);
	alias XbG_H0 : voltage is Vneg_temp(0);
	alias XbG_H1 : voltage is Vneg_temp(1);
	alias XbG_H2 : voltage is Vneg_temp(2);
	alias XbG_H3 : voltage is Vneg_temp(3);
	alias XbG_H4 : voltage is Vneg_temp(4);
	alias XbG_H5 : voltage is Vneg_temp(5);
	alias XbG_H6 : voltage is Vneg_temp(6);
	alias XbG_H7 : voltage is Vneg_temp(7);
	alias XbG_H8 : voltage is Vneg_temp(8);
	alias XbG_H9 : voltage is Vneg_temp(9);
	alias XbG_H10 : voltage is Vneg_temp(10);
	alias XbG_H11 : voltage is Vneg_temp(11);
	alias XbG_H12 : voltage is Vneg_temp(12);
	alias XbG_H13 : voltage is Vneg_temp(13);
	alias XbG_H14 : voltage is Vneg_temp(14);
	alias XbG_H15 : voltage is Vneg_temp(15);
	alias XbG_H16 : voltage is Vneg_temp(16);
	alias XbG_H17 : voltage is Vneg_temp(17);
	alias XbG_H18 : voltage is Vneg_temp(18);
	alias XbG_H19 : voltage is Vneg_temp(19);
	alias XbG_H20 : voltage is Vneg_temp(20);
	alias XbG_H21 : voltage is Vneg_temp(21);
	alias XbG_H22 : voltage is Vneg_temp(22);
	alias XbG_H23 : voltage is Vneg_temp(23);
	alias XbG_H24 : voltage is Vneg_temp(24);
	alias XbG_H25 : voltage is Vneg_temp(25);
	alias XbG_H26 : voltage is Vneg_temp(26);
	alias XbG_H27 : voltage is Vneg_temp(27);
	alias XbG_H28 : voltage is Vneg_temp(28);
	alias XbG_H29 : voltage is Vneg_temp(29);
	alias XbG_H30 : voltage is Vneg_temp(30);
	alias XbG_H31 : voltage is Vneg_temp(31);
	alias XbG_H32 : voltage is Vneg_temp(32);
	alias XbG_H33 : voltage is Vneg_temp(33);
	alias XbG_H34 : voltage is Vneg_temp(34);
	alias XbG_H35 : voltage is Vneg_temp(35);
	alias XbG_H36 : voltage is Vneg_temp(36);
	alias XbG_H37 : voltage is Vneg_temp(37);
	alias XbG_H38 : voltage is Vneg_temp(38);
	alias XbG_H39 : voltage is Vneg_temp(39);
	alias XbG_H40 : voltage is Vneg_temp(40);
	alias XbG_H41 : voltage is Vneg_temp(41);
	alias XbG_H42 : voltage is Vneg_temp(42);
	alias XbG_H43 : voltage is Vneg_temp(43);
	alias XbG_H44 : voltage is Vneg_temp(44);
	alias XbG_H45 : voltage is Vneg_temp(45);
	alias XbG_H46 : voltage is Vneg_temp(46);
	alias XbG_H47 : voltage is Vneg_temp(47);
	alias XbG_H48 : voltage is Vneg_temp(48);
	alias XbG_H49 : voltage is Vneg_temp(49);
	alias XbG_H50 : voltage is Vneg_temp(50);
	alias XbG_H51 : voltage is Vneg_temp(51);
	alias XbG_H52 : voltage is Vneg_temp(52);
	alias XbG_H53 : voltage is Vneg_temp(53);
	alias XbG_H54 : voltage is Vneg_temp(54);
	alias XbG_H55 : voltage is Vneg_temp(55);
	alias XbG_H56 : voltage is Vneg_temp(56);
	alias XbG_H57 : voltage is Vneg_temp(57);
	alias XbG_H58 : voltage is Vneg_temp(58);
	alias XbG_H59 : voltage is Vneg_temp(59);
	alias XbG_H60 : voltage is Vneg_temp(60);
	alias XbG_H61 : voltage is Vneg_temp(61);
	alias XbG_H62 : voltage is Vneg_temp(62);
	alias XbG_H63 : voltage is Vneg_temp(63);
	alias XbG_H64 : voltage is Vneg_temp(64);
	alias XbG_H65 : voltage is Vneg_temp(65);
	alias XbG_H66 : voltage is Vneg_temp(66);
	alias XbG_H67 : voltage is Vneg_temp(67);
	alias XbG_H68 : voltage is Vneg_temp(68);
	alias XbG_H69 : voltage is Vneg_temp(69);
	alias XbG_H70 : voltage is Vneg_temp(70);
	alias XbG_H71 : voltage is Vneg_temp(71);
	alias XbG_H72 : voltage is Vneg_temp(72);
	alias XbG_H73 : voltage is Vneg_temp(73);
	alias XbG_H74 : voltage is Vneg_temp(74);
	alias XbG_H75 : voltage is Vneg_temp(75);
	alias XbG_H76 : voltage is Vneg_temp(76);
	alias XbG_H77 : voltage is Vneg_temp(77);
	alias XbG_H78 : voltage is Vneg_temp(78);
	alias XbG_H79 : voltage is Vneg_temp(79);
	alias XbG_H80 : voltage is Vneg_temp(80);
	alias XbG_H81 : voltage is Vneg_temp(81);
	alias XbG_H82 : voltage is Vneg_temp(82);
	alias XbG_H83 : voltage is Vneg_temp(83);
	alias XbG_H84 : voltage is Vneg_temp(84);
	alias XbG_H85 : voltage is Vneg_temp(85);
	alias XbG_H86 : voltage is Vneg_temp(86);
	alias XbG_H87 : voltage is Vneg_temp(87);
	alias XbG_H88 : voltage is Vneg_temp(88);
	alias XbG_H89 : voltage is Vneg_temp(89);
	alias XbG_H90 : voltage is Vneg_temp(90);
	alias XbG_H91 : voltage is Vneg_temp(91);
	alias XbG_H92 : voltage is Vneg_temp(92);
	alias XbG_H93 : voltage is Vneg_temp(93);
	alias XbG_H94 : voltage is Vneg_temp(94);
	alias XbG_H95 : voltage is Vneg_temp(95);
	alias XbG_H96 : voltage is Vneg_temp(96);
	alias XbG_H97 : voltage is Vneg_temp(97);
	alias XbG_H98 : voltage is Vneg_temp(98);
	alias XbG_H99 : voltage is Vneg_temp(99);
	alias XbG_H100 : voltage is Vneg_temp(100);
	alias XbG_H101 : voltage is Vneg_temp(101);
	alias XbG_H102 : voltage is Vneg_temp(102);
	alias XbG_H103 : voltage is Vneg_temp(103);
	alias XbG_H104 : voltage is Vneg_temp(104);
	alias XbG_H105 : voltage is Vneg_temp(105);
	alias XbG_H106 : voltage is Vneg_temp(106);
	alias XbG_H107 : voltage is Vneg_temp(107);
	alias XbG_H108 : voltage is Vneg_temp(108);
	alias XbG_H109 : voltage is Vneg_temp(109);
	alias XbG_H110 : voltage is Vneg_temp(110);
	alias XbG_H111 : voltage is Vneg_temp(111);
	alias XbG_H112 : voltage is Vneg_temp(112);
	alias XbG_H113 : voltage is Vneg_temp(113);
	alias XbG_H114 : voltage is Vneg_temp(114);
	alias XbG_H115 : voltage is Vneg_temp(115);
	alias XbG_H116 : voltage is Vneg_temp(116);
	alias XbG_H117 : voltage is Vneg_temp(117);
	alias XbG_H118 : voltage is Vneg_temp(118);
	alias XbG_H119 : voltage is Vneg_temp(119);
	alias XbG_H120 : voltage is Vneg_temp(120);
	alias XbG_H121 : voltage is Vneg_temp(121);
	alias XbG_H122 : voltage is Vneg_temp(122);
	alias XbG_H123 : voltage is Vneg_temp(123);
	alias XbG_H124 : voltage is Vneg_temp(124);
	alias XbG_H125 : voltage is Vneg_temp(125);
	alias XbG_H126 : voltage is Vneg_temp(126);
	alias XbG_H127 : voltage is Vneg_temp(127);
	alias XbG_H128 : voltage is Vneg_temp(128);
	alias XbG_H129 : voltage is Vneg_temp(129);
	alias XbG_H130 : voltage is Vneg_temp(130);
	alias XbG_H131 : voltage is Vneg_temp(131);
	alias XbG_H132 : voltage is Vneg_temp(132);
	alias XbG_H133 : voltage is Vneg_temp(133);
	alias XbG_H134 : voltage is Vneg_temp(134);
	alias XbG_H135 : voltage is Vneg_temp(135);
	alias XbG_H136 : voltage is Vneg_temp(136);
	alias XbG_H137 : voltage is Vneg_temp(137);
	alias XbG_H138 : voltage is Vneg_temp(138);
	alias XbG_H139 : voltage is Vneg_temp(139);
	alias XbG_H140 : voltage is Vneg_temp(140);
	alias XbG_H141 : voltage is Vneg_temp(141);
	alias XbG_H142 : voltage is Vneg_temp(142);
	alias XbG_H143 : voltage is Vneg_temp(143);
	alias XbG_H144 : voltage is Vneg_temp(144);
	alias XbG_H145 : voltage is Vneg_temp(145);
	alias XbG_H146 : voltage is Vneg_temp(146);
	alias XbG_H147 : voltage is Vneg_temp(147);
	alias XbG_H148 : voltage is Vneg_temp(148);
	alias XbG_H149 : voltage is Vneg_temp(149);
	alias XbG_H150 : voltage is Vneg_temp(150);
	alias XbG_H151 : voltage is Vneg_temp(151);
	alias XbG_H152 : voltage is Vneg_temp(152);
	alias XbG_H153 : voltage is Vneg_temp(153);
	alias XbG_H154 : voltage is Vneg_temp(154);
	alias XbG_H155 : voltage is Vneg_temp(155);
	alias XbG_H156 : voltage is Vneg_temp(156);
	alias XbG_H157 : voltage is Vneg_temp(157);
	alias XbG_H158 : voltage is Vneg_temp(158);
	alias XbG_H159 : voltage is Vneg_temp(159);
	alias XbG_H160 : voltage is Vneg_temp(160);
	alias XbG_H161 : voltage is Vneg_temp(161);
	alias XbG_H162 : voltage is Vneg_temp(162);
	alias XbG_H163 : voltage is Vneg_temp(163);
	alias XbG_H164 : voltage is Vneg_temp(164);
	alias XbG_H165 : voltage is Vneg_temp(165);
	alias XbG_H166 : voltage is Vneg_temp(166);
	alias XbG_H167 : voltage is Vneg_temp(167);
	alias XbG_H168 : voltage is Vneg_temp(168);
	alias XbG_H169 : voltage is Vneg_temp(169);
	alias XbG_H170 : voltage is Vneg_temp(170);
	alias XbG_H171 : voltage is Vneg_temp(171);
	alias XbG_H172 : voltage is Vneg_temp(172);
	alias XbG_H173 : voltage is Vneg_temp(173);
	alias XbG_H174 : voltage is Vneg_temp(174);
	alias XbG_H175 : voltage is Vneg_temp(175);
	alias XbG_H176 : voltage is Vneg_temp(176);
	alias XbG_H177 : voltage is Vneg_temp(177);
	alias XbG_H178 : voltage is Vneg_temp(178);
	alias XbG_H179 : voltage is Vneg_temp(179);
	alias XbG_H180 : voltage is Vneg_temp(180);
	alias XbG_H181 : voltage is Vneg_temp(181);
	alias XbG_H182 : voltage is Vneg_temp(182);
	alias XbG_H183 : voltage is Vneg_temp(183);
	alias XbG_H184 : voltage is Vneg_temp(184);
	alias XbG_H185 : voltage is Vneg_temp(185);
	alias XbG_H186 : voltage is Vneg_temp(186);
	alias XbG_H187 : voltage is Vneg_temp(187);
	alias XbG_H188 : voltage is Vneg_temp(188);
	alias XbG_H189 : voltage is Vneg_temp(189);
	alias XbG_H190 : voltage is Vneg_temp(190);
	alias XbG_H191 : voltage is Vneg_temp(191);
	alias XbG_H192 : voltage is Vneg_temp(192);
	alias XbG_H193 : voltage is Vneg_temp(193);
	alias XbG_H194 : voltage is Vneg_temp(194);
	alias XbG_H195 : voltage is Vneg_temp(195);
	alias XbG_H196 : voltage is Vneg_temp(196);
	alias XbG_H197 : voltage is Vneg_temp(197);
	alias XbG_H198 : voltage is Vneg_temp(198);
	alias XbG_H199 : voltage is Vneg_temp(199);
	alias XbG_H200 : voltage is Vneg_temp(200);
	alias XbG_H201 : voltage is Vneg_temp(201);
	alias XbG_H202 : voltage is Vneg_temp(202);
	alias XbG_H203 : voltage is Vneg_temp(203);
	alias XbG_H204 : voltage is Vneg_temp(204);
	alias XbG_H205 : voltage is Vneg_temp(205);
	alias XbG_H206 : voltage is Vneg_temp(206);
	alias XbG_H207 : voltage is Vneg_temp(207);
	alias XbG_H208 : voltage is Vneg_temp(208);
	alias XbG_H209 : voltage is Vneg_temp(209);
	alias XbG_H210 : voltage is Vneg_temp(210);
	alias XbG_H211 : voltage is Vneg_temp(211);
	alias XbG_H212 : voltage is Vneg_temp(212);
	alias XbG_H213 : voltage is Vneg_temp(213);
	alias XbG_H214 : voltage is Vneg_temp(214);
	alias XbG_H215 : voltage is Vneg_temp(215);
	alias XbG_H216 : voltage is Vneg_temp(216);
	alias XbG_H217 : voltage is Vneg_temp(217);
	alias XbG_H218 : voltage is Vneg_temp(218);
	alias XbG_H219 : voltage is Vneg_temp(219);
	alias XbG_H220 : voltage is Vneg_temp(220);
	alias XbG_H221 : voltage is Vneg_temp(221);
	alias XbG_H222 : voltage is Vneg_temp(222);
	alias XbG_H223 : voltage is Vneg_temp(223);
	alias XbG_H224 : voltage is Vneg_temp(224);
	alias XbG_H225 : voltage is Vneg_temp(225);
	alias XbG_H226 : voltage is Vneg_temp(226);
	alias XbG_H227 : voltage is Vneg_temp(227);
	alias XbG_H228 : voltage is Vneg_temp(228);
	alias XbG_H229 : voltage is Vneg_temp(229);
	alias XbG_H230 : voltage is Vneg_temp(230);
	alias XbG_H231 : voltage is Vneg_temp(231);
	alias XbG_H232 : voltage is Vneg_temp(232);
	alias XbG_H233 : voltage is Vneg_temp(233);
	alias XbG_H234 : voltage is Vneg_temp(234);
	alias XbG_H235 : voltage is Vneg_temp(235);
	alias XbG_H236 : voltage is Vneg_temp(236);
	alias XbG_H237 : voltage is Vneg_temp(237);
	alias XbG_H238 : voltage is Vneg_temp(238);
	alias XbG_H239 : voltage is Vneg_temp(239);
	alias XbG_H240 : voltage is Vneg_temp(240);
	alias XbG_H241 : voltage is Vneg_temp(241);
	alias XbG_H242 : voltage is Vneg_temp(242);
	alias XbG_H243 : voltage is Vneg_temp(243);
	alias XbG_H244 : voltage is Vneg_temp(244);
	alias XbG_H245 : voltage is Vneg_temp(245);
	alias XbG_H246 : voltage is Vneg_temp(246);
	alias XbG_H247 : voltage is Vneg_temp(247);
	alias XbG_H248 : voltage is Vneg_temp(248);
	alias XbG_H249 : voltage is Vneg_temp(249);
	alias XbG_H250 : voltage is Vneg_temp(250);
	alias XbG_H251 : voltage is Vneg_temp(251);
	alias XbG_H252 : voltage is Vneg_temp(252);
	alias XbG_H253 : voltage is Vneg_temp(253);
	alias XbG_H254 : voltage is Vneg_temp(254);
	alias XbG_H255 : voltage is Vneg_temp(255);
	alias XbG_H256 : voltage is Vneg_temp(256);
	alias XbG_H257 : voltage is Vneg_temp(257);
	alias XbG_H258 : voltage is Vneg_temp(258);
	alias XbG_H259 : voltage is Vneg_temp(259);
	alias XbG_H260 : voltage is Vneg_temp(260);
	alias XbG_H261 : voltage is Vneg_temp(261);
	alias XbG_H262 : voltage is Vneg_temp(262);
	alias XbG_H263 : voltage is Vneg_temp(263);
	alias XbG_H264 : voltage is Vneg_temp(264);
	alias XbG_H265 : voltage is Vneg_temp(265);
	alias XbG_H266 : voltage is Vneg_temp(266);
	alias XbG_H267 : voltage is Vneg_temp(267);
	alias XbG_H268 : voltage is Vneg_temp(268);
	alias XbG_H269 : voltage is Vneg_temp(269);
	alias XbG_H270 : voltage is Vneg_temp(270);
	alias XbG_H271 : voltage is Vneg_temp(271);
	alias XbG_H272 : voltage is Vneg_temp(272);
	alias XbG_H273 : voltage is Vneg_temp(273);
	alias XbG_H274 : voltage is Vneg_temp(274);
	alias XbG_H275 : voltage is Vneg_temp(275);
	alias XbG_H276 : voltage is Vneg_temp(276);
	alias XbG_H277 : voltage is Vneg_temp(277);
	alias XbG_H278 : voltage is Vneg_temp(278);
	alias XbG_H279 : voltage is Vneg_temp(279);
	alias XbG_H280 : voltage is Vneg_temp(280);
	alias XbG_H281 : voltage is Vneg_temp(281);
	alias XbG_H282 : voltage is Vneg_temp(282);
	alias XbG_H283 : voltage is Vneg_temp(283);
	alias XbG_H284 : voltage is Vneg_temp(284);
	alias XbG_H285 : voltage is Vneg_temp(285);
	alias XbG_H286 : voltage is Vneg_temp(286);
	alias XbG_H287 : voltage is Vneg_temp(287);
	alias XbG_H288 : voltage is Vneg_temp(288);
	alias XbG_H289 : voltage is Vneg_temp(289);
	alias XbG_H290 : voltage is Vneg_temp(290);
	alias XbG_H291 : voltage is Vneg_temp(291);
	alias XbG_H292 : voltage is Vneg_temp(292);
	alias XbG_H293 : voltage is Vneg_temp(293);
	alias XbG_H294 : voltage is Vneg_temp(294);
	alias XbG_H295 : voltage is Vneg_temp(295);
	alias XbG_H296 : voltage is Vneg_temp(296);
	alias XbG_H297 : voltage is Vneg_temp(297);
	alias XbG_H298 : voltage is Vneg_temp(298);
	alias XbG_H299 : voltage is Vneg_temp(299);
	alias XbG_H300 : voltage is Vneg_temp(300);
	alias XbG_H301 : voltage is Vneg_temp(301);
	alias XbG_H302 : voltage is Vneg_temp(302);
	alias XbG_H303 : voltage is Vneg_temp(303);
	alias XbG_H304 : voltage is Vneg_temp(304);
	alias XbG_H305 : voltage is Vneg_temp(305);
	alias XbG_H306 : voltage is Vneg_temp(306);
	alias XbG_H307 : voltage is Vneg_temp(307);
	alias XbG_H308 : voltage is Vneg_temp(308);
	alias XbG_H309 : voltage is Vneg_temp(309);
	alias XbG_H310 : voltage is Vneg_temp(310);
	alias XbG_H311 : voltage is Vneg_temp(311);
	alias XbG_H312 : voltage is Vneg_temp(312);
	alias XbG_H313 : voltage is Vneg_temp(313);
	alias XbG_H314 : voltage is Vneg_temp(314);
	alias XbG_H315 : voltage is Vneg_temp(315);
	alias XbG_H316 : voltage is Vneg_temp(316);
	alias XbG_H317 : voltage is Vneg_temp(317);
	alias XbG_H318 : voltage is Vneg_temp(318);
	alias XbG_H319 : voltage is Vneg_temp(319);
	alias XbG_H320 : voltage is Vneg_temp(320);
	alias XbG_H321 : voltage is Vneg_temp(321);
	alias XbG_H322 : voltage is Vneg_temp(322);
	alias XbG_H323 : voltage is Vneg_temp(323);
	alias XbG_H324 : voltage is Vneg_temp(324);
	alias XbG_H325 : voltage is Vneg_temp(325);
	alias XbG_H326 : voltage is Vneg_temp(326);
	alias XbG_H327 : voltage is Vneg_temp(327);
	alias XbG_H328 : voltage is Vneg_temp(328);
	alias XbG_H329 : voltage is Vneg_temp(329);
	alias XbG_H330 : voltage is Vneg_temp(330);
	alias XbG_H331 : voltage is Vneg_temp(331);
	alias XbG_H332 : voltage is Vneg_temp(332);
	alias XbG_H333 : voltage is Vneg_temp(333);
	alias XbG_H334 : voltage is Vneg_temp(334);
	alias XbG_H335 : voltage is Vneg_temp(335);
	alias XbG_H336 : voltage is Vneg_temp(336);
	alias XbG_H337 : voltage is Vneg_temp(337);
	alias XbG_H338 : voltage is Vneg_temp(338);
	alias XbG_H339 : voltage is Vneg_temp(339);
	alias XbG_H340 : voltage is Vneg_temp(340);
	alias XbG_H341 : voltage is Vneg_temp(341);
	alias XbG_H342 : voltage is Vneg_temp(342);
	alias XbG_H343 : voltage is Vneg_temp(343);
	alias XbG_H344 : voltage is Vneg_temp(344);
	alias XbG_H345 : voltage is Vneg_temp(345);
	alias XbG_H346 : voltage is Vneg_temp(346);
	alias XbG_H347 : voltage is Vneg_temp(347);
	alias XbG_H348 : voltage is Vneg_temp(348);
	alias XbG_H349 : voltage is Vneg_temp(349);
	alias XbG_H350 : voltage is Vneg_temp(350);
	alias XbG_H351 : voltage is Vneg_temp(351);
	alias XbG_H352 : voltage is Vneg_temp(352);
	alias XbG_H353 : voltage is Vneg_temp(353);
	alias XbG_H354 : voltage is Vneg_temp(354);
	alias XbG_H355 : voltage is Vneg_temp(355);
	alias XbG_H356 : voltage is Vneg_temp(356);
	alias XbG_H357 : voltage is Vneg_temp(357);
	alias XbG_H358 : voltage is Vneg_temp(358);
	alias XbG_H359 : voltage is Vneg_temp(359);
	alias XbG_H360 : voltage is Vneg_temp(360);
	alias XbG_H361 : voltage is Vneg_temp(361);
	alias XbG_H362 : voltage is Vneg_temp(362);
	alias XbG_H363 : voltage is Vneg_temp(363);
	alias XbG_H364 : voltage is Vneg_temp(364);
	alias XbG_H365 : voltage is Vneg_temp(365);
	alias XbG_H366 : voltage is Vneg_temp(366);
	alias XbG_H367 : voltage is Vneg_temp(367);
	alias XbG_H368 : voltage is Vneg_temp(368);
	alias XbG_H369 : voltage is Vneg_temp(369);
	alias XbG_H370 : voltage is Vneg_temp(370);
	alias XbG_H371 : voltage is Vneg_temp(371);
	alias XbG_H372 : voltage is Vneg_temp(372);
	alias XbG_H373 : voltage is Vneg_temp(373);
	alias XbG_H374 : voltage is Vneg_temp(374);
	alias XbG_H375 : voltage is Vneg_temp(375);
	alias XbG_H376 : voltage is Vneg_temp(376);
	alias XbG_H377 : voltage is Vneg_temp(377);
	alias XbG_H378 : voltage is Vneg_temp(378);
	alias XbG_H379 : voltage is Vneg_temp(379);
	alias XbG_H380 : voltage is Vneg_temp(380);
	alias XbG_H381 : voltage is Vneg_temp(381);
	alias XbG_H382 : voltage is Vneg_temp(382);
	alias XbG_H383 : voltage is Vneg_temp(383);
	alias XbG_H384 : voltage is Vneg_temp(384);
	alias XbG_H385 : voltage is Vneg_temp(385);
	alias XbG_H386 : voltage is Vneg_temp(386);
	alias XbG_H387 : voltage is Vneg_temp(387);
	alias XbG_H388 : voltage is Vneg_temp(388);
	alias XbG_H389 : voltage is Vneg_temp(389);
	alias XbG_H390 : voltage is Vneg_temp(390);
	alias XbG_H391 : voltage is Vneg_temp(391);
	alias XbG_H392 : voltage is Vneg_temp(392);
	alias XbG_H393 : voltage is Vneg_temp(393);
	alias XbG_H394 : voltage is Vneg_temp(394);
	alias XbG_H395 : voltage is Vneg_temp(395);
	alias XbG_H396 : voltage is Vneg_temp(396);
	alias XbG_H397 : voltage is Vneg_temp(397);
	alias XbG_H398 : voltage is Vneg_temp(398);
	alias XbG_H399 : voltage is Vneg_temp(399);
	alias XbG_H400 : voltage is Vneg_temp(400);
	alias XbG_H401 : voltage is Vneg_temp(401);
	alias XbG_H402 : voltage is Vneg_temp(402);
	alias XbG_H403 : voltage is Vneg_temp(403);
	alias XbG_H404 : voltage is Vneg_temp(404);
	alias XbG_H405 : voltage is Vneg_temp(405);
	alias XbG_H406 : voltage is Vneg_temp(406);
	alias XbG_H407 : voltage is Vneg_temp(407);
	alias XbG_H408 : voltage is Vneg_temp(408);
	alias XbG_H409 : voltage is Vneg_temp(409);
	alias XbG_H410 : voltage is Vneg_temp(410);
	alias XbG_H411 : voltage is Vneg_temp(411);
	alias XbG_H412 : voltage is Vneg_temp(412);
	alias XbG_H413 : voltage is Vneg_temp(413);
	alias XbG_H414 : voltage is Vneg_temp(414);
	alias XbG_H415 : voltage is Vneg_temp(415);
	alias XbG_H416 : voltage is Vneg_temp(416);
	alias XbG_H417 : voltage is Vneg_temp(417);
	alias XbG_H418 : voltage is Vneg_temp(418);
	alias XbG_H419 : voltage is Vneg_temp(419);
	alias XbG_H420 : voltage is Vneg_temp(420);
	alias XbG_H421 : voltage is Vneg_temp(421);
	alias XbG_H422 : voltage is Vneg_temp(422);
	alias XbG_H423 : voltage is Vneg_temp(423);
	alias XbG_H424 : voltage is Vneg_temp(424);
	alias XbG_H425 : voltage is Vneg_temp(425);
	alias XbG_H426 : voltage is Vneg_temp(426);
	alias XbG_H427 : voltage is Vneg_temp(427);
	alias XbG_H428 : voltage is Vneg_temp(428);
	alias XbG_H429 : voltage is Vneg_temp(429);
	alias XbG_H430 : voltage is Vneg_temp(430);
	alias XbG_H431 : voltage is Vneg_temp(431);
	alias XbG_H432 : voltage is Vneg_temp(432);
	alias XbG_H433 : voltage is Vneg_temp(433);
	alias XbG_H434 : voltage is Vneg_temp(434);
	alias XbG_H435 : voltage is Vneg_temp(435);
	alias XbG_H436 : voltage is Vneg_temp(436);
	alias XbG_H437 : voltage is Vneg_temp(437);
	alias XbG_H438 : voltage is Vneg_temp(438);
	alias XbG_H439 : voltage is Vneg_temp(439);
	alias XbG_H440 : voltage is Vneg_temp(440);
	alias XbG_H441 : voltage is Vneg_temp(441);
	alias XbG_H442 : voltage is Vneg_temp(442);
	alias XbG_H443 : voltage is Vneg_temp(443);
	alias XbG_H444 : voltage is Vneg_temp(444);
	alias XbG_H445 : voltage is Vneg_temp(445);
	alias XbG_H446 : voltage is Vneg_temp(446);
	alias XbG_H447 : voltage is Vneg_temp(447);
	alias XbG_H448 : voltage is Vneg_temp(448);
	alias XbG_H449 : voltage is Vneg_temp(449);
	alias XbG_H450 : voltage is Vneg_temp(450);
	alias XbG_H451 : voltage is Vneg_temp(451);
	alias XbG_H452 : voltage is Vneg_temp(452);
	alias XbG_H453 : voltage is Vneg_temp(453);
	alias XbG_H454 : voltage is Vneg_temp(454);
	alias XbG_H455 : voltage is Vneg_temp(455);
	alias XbG_H456 : voltage is Vneg_temp(456);
	alias XbG_H457 : voltage is Vneg_temp(457);
	alias XbG_H458 : voltage is Vneg_temp(458);
	alias XbG_H459 : voltage is Vneg_temp(459);
	alias XbG_H460 : voltage is Vneg_temp(460);
	alias XbG_H461 : voltage is Vneg_temp(461);
	alias XbG_H462 : voltage is Vneg_temp(462);
	alias XbG_H463 : voltage is Vneg_temp(463);
	alias XbG_H464 : voltage is Vneg_temp(464);
	alias XbG_H465 : voltage is Vneg_temp(465);
	alias XbG_H466 : voltage is Vneg_temp(466);
	alias XbG_H467 : voltage is Vneg_temp(467);
	alias XbG_H468 : voltage is Vneg_temp(468);
	alias XbG_H469 : voltage is Vneg_temp(469);
	alias XbG_H470 : voltage is Vneg_temp(470);
	alias XbG_H471 : voltage is Vneg_temp(471);
	alias XbG_H472 : voltage is Vneg_temp(472);
	alias XbG_H473 : voltage is Vneg_temp(473);
	alias XbG_H474 : voltage is Vneg_temp(474);
	alias XbG_H475 : voltage is Vneg_temp(475);
	alias XbG_H476 : voltage is Vneg_temp(476);
	alias XbG_H477 : voltage is Vneg_temp(477);
	alias XbG_H478 : voltage is Vneg_temp(478);
	alias XbG_H479 : voltage is Vneg_temp(479);
	alias XbG_H480 : voltage is Vneg_temp(480);
	alias XbG_H481 : voltage is Vneg_temp(481);
	alias XbG_H482 : voltage is Vneg_temp(482);
	alias XbG_H483 : voltage is Vneg_temp(483);
	alias XbG_H484 : voltage is Vneg_temp(484);
	alias XbG_H485 : voltage is Vneg_temp(485);
	alias XbG_H486 : voltage is Vneg_temp(486);
	alias XbG_H487 : voltage is Vneg_temp(487);
	alias XbG_H488 : voltage is Vneg_temp(488);
	alias XbG_H489 : voltage is Vneg_temp(489);
	alias XbG_H490 : voltage is Vneg_temp(490);
	alias XbG_H491 : voltage is Vneg_temp(491);
	alias XbG_H492 : voltage is Vneg_temp(492);
	alias XbG_H493 : voltage is Vneg_temp(493);
	alias XbG_H494 : voltage is Vneg_temp(494);
	alias XbG_H495 : voltage is Vneg_temp(495);
	alias XbG_H496 : voltage is Vneg_temp(496);
	alias XbG_H497 : voltage is Vneg_temp(497);
	alias XbG_H498 : voltage is Vneg_temp(498);
	alias XbG_H499 : voltage is Vneg_temp(499);
	alias XbG_H500 : voltage is Vneg_temp(500);
	alias XbG_H501 : voltage is Vneg_temp(501);
	alias XbG_H502 : voltage is Vneg_temp(502);
	alias XbG_H503 : voltage is Vneg_temp(503);
	alias XbG_H504 : voltage is Vneg_temp(504);
	alias XbG_H505 : voltage is Vneg_temp(505);
	alias XbG_H506 : voltage is Vneg_temp(506);
	alias XbG_H507 : voltage is Vneg_temp(507);
	alias XbG_H508 : voltage is Vneg_temp(508);
	alias XbG_H509 : voltage is Vneg_temp(509);
	alias XbG_H510 : voltage is Vneg_temp(510);
	alias XbG_H511 : voltage is Vneg_temp(511);
	alias XbG_H512 : voltage is Vneg_temp(512);
	alias XbG_H513 : voltage is Vneg_temp(513);
	alias XbG_H514 : voltage is Vneg_temp(514);
	alias XbG_H515 : voltage is Vneg_temp(515);
	alias XbG_H516 : voltage is Vneg_temp(516);
	alias XbG_H517 : voltage is Vneg_temp(517);
	alias XbG_H518 : voltage is Vneg_temp(518);
	alias XbG_H519 : voltage is Vneg_temp(519);
	alias XbG_H520 : voltage is Vneg_temp(520);
	alias XbG_H521 : voltage is Vneg_temp(521);
	alias XbG_H522 : voltage is Vneg_temp(522);
	alias XbG_H523 : voltage is Vneg_temp(523);
	alias XbG_H524 : voltage is Vneg_temp(524);
	alias XbG_H525 : voltage is Vneg_temp(525);
	alias XbG_H526 : voltage is Vneg_temp(526);
	alias XbG_H527 : voltage is Vneg_temp(527);
	alias XbG_H528 : voltage is Vneg_temp(528);
	alias XbG_H529 : voltage is Vneg_temp(529);
	alias XbG_H530 : voltage is Vneg_temp(530);
	alias XbG_H531 : voltage is Vneg_temp(531);
	alias XbG_H532 : voltage is Vneg_temp(532);
	alias XbG_H533 : voltage is Vneg_temp(533);
	alias XbG_H534 : voltage is Vneg_temp(534);
	alias XbG_H535 : voltage is Vneg_temp(535);
	alias XbG_H536 : voltage is Vneg_temp(536);
	alias XbG_H537 : voltage is Vneg_temp(537);
	alias XbG_H538 : voltage is Vneg_temp(538);
	alias XbG_H539 : voltage is Vneg_temp(539);
	alias XbG_H540 : voltage is Vneg_temp(540);
	alias XbG_H541 : voltage is Vneg_temp(541);
	alias XbG_H542 : voltage is Vneg_temp(542);
	alias XbG_H543 : voltage is Vneg_temp(543);
	alias XbG_H544 : voltage is Vneg_temp(544);
	alias XbG_H545 : voltage is Vneg_temp(545);
	alias XbG_H546 : voltage is Vneg_temp(546);
	alias XbG_H547 : voltage is Vneg_temp(547);
	alias XbG_H548 : voltage is Vneg_temp(548);
	alias XbG_H549 : voltage is Vneg_temp(549);
	alias XbG_H550 : voltage is Vneg_temp(550);
	alias XbG_H551 : voltage is Vneg_temp(551);
	alias XbG_H552 : voltage is Vneg_temp(552);
	alias XbG_H553 : voltage is Vneg_temp(553);
	alias XbG_H554 : voltage is Vneg_temp(554);
	alias XbG_H555 : voltage is Vneg_temp(555);
	alias XbG_H556 : voltage is Vneg_temp(556);
	alias XbG_H557 : voltage is Vneg_temp(557);
	alias XbG_H558 : voltage is Vneg_temp(558);
	alias XbG_H559 : voltage is Vneg_temp(559);
	alias XbG_H560 : voltage is Vneg_temp(560);
	alias XbG_H561 : voltage is Vneg_temp(561);
	alias XbG_H562 : voltage is Vneg_temp(562);
	alias XbG_H563 : voltage is Vneg_temp(563);
	alias XbG_H564 : voltage is Vneg_temp(564);
	alias XbG_H565 : voltage is Vneg_temp(565);
	alias XbG_H566 : voltage is Vneg_temp(566);
	alias XbG_H567 : voltage is Vneg_temp(567);
	alias XbG_H568 : voltage is Vneg_temp(568);
	alias XbG_H569 : voltage is Vneg_temp(569);
	alias XbG_H570 : voltage is Vneg_temp(570);
	alias XbG_H571 : voltage is Vneg_temp(571);
	alias XbG_H572 : voltage is Vneg_temp(572);
	alias XbG_H573 : voltage is Vneg_temp(573);
	alias XbG_H574 : voltage is Vneg_temp(574);
	alias XbG_H575 : voltage is Vneg_temp(575);
	alias XbG_H576 : voltage is Vneg_temp(576);
	alias XbG_H577 : voltage is Vneg_temp(577);
	alias XbG_H578 : voltage is Vneg_temp(578);
	alias XbG_H579 : voltage is Vneg_temp(579);
	alias XbG_H580 : voltage is Vneg_temp(580);
	alias XbG_H581 : voltage is Vneg_temp(581);
	alias XbG_H582 : voltage is Vneg_temp(582);
	alias XbG_H583 : voltage is Vneg_temp(583);
	alias XbG_H584 : voltage is Vneg_temp(584);
	alias XbG_H585 : voltage is Vneg_temp(585);
	alias XbG_H586 : voltage is Vneg_temp(586);
	alias XbG_H587 : voltage is Vneg_temp(587);
	alias XbG_H588 : voltage is Vneg_temp(588);
	alias XbG_H589 : voltage is Vneg_temp(589);
	alias XbG_H590 : voltage is Vneg_temp(590);
	alias XbG_H591 : voltage is Vneg_temp(591);
	alias XbG_H592 : voltage is Vneg_temp(592);
	alias XbG_H593 : voltage is Vneg_temp(593);
	alias XbG_H594 : voltage is Vneg_temp(594);
	alias XbG_H595 : voltage is Vneg_temp(595);
	alias XbG_H596 : voltage is Vneg_temp(596);
	alias XbG_H597 : voltage is Vneg_temp(597);
	alias XbG_H598 : voltage is Vneg_temp(598);
	alias XbG_H599 : voltage is Vneg_temp(599);
	alias XbG_H600 : voltage is Vneg_temp(600);
	alias XbG_H601 : voltage is Vneg_temp(601);
	alias XbG_H602 : voltage is Vneg_temp(602);
	alias XbG_H603 : voltage is Vneg_temp(603);
	alias XbG_H604 : voltage is Vneg_temp(604);
	alias XbG_H605 : voltage is Vneg_temp(605);
	alias XbG_H606 : voltage is Vneg_temp(606);
	alias XbG_H607 : voltage is Vneg_temp(607);
	alias XbG_H608 : voltage is Vneg_temp(608);
	alias XbG_H609 : voltage is Vneg_temp(609);
	alias XbG_H610 : voltage is Vneg_temp(610);
	alias XbG_H611 : voltage is Vneg_temp(611);
	alias XbG_H612 : voltage is Vneg_temp(612);
	alias XbG_H613 : voltage is Vneg_temp(613);
	alias XbG_H614 : voltage is Vneg_temp(614);
	alias XbG_H615 : voltage is Vneg_temp(615);
	alias XbG_H616 : voltage is Vneg_temp(616);
	alias XbG_H617 : voltage is Vneg_temp(617);
	alias XbG_H618 : voltage is Vneg_temp(618);
	alias XbG_H619 : voltage is Vneg_temp(619);
	alias XbG_H620 : voltage is Vneg_temp(620);
	alias XbG_H621 : voltage is Vneg_temp(621);
	alias XbG_H622 : voltage is Vneg_temp(622);
	alias XbG_H623 : voltage is Vneg_temp(623);
	alias XbG_H624 : voltage is Vneg_temp(624);
	alias XbG_H625 : voltage is Vneg_temp(625);
	alias XbG_H626 : voltage is Vneg_temp(626);
	alias XbG_H627 : voltage is Vneg_temp(627);
	alias XbG_H628 : voltage is Vneg_temp(628);
	alias XbG_H629 : voltage is Vneg_temp(629);
	alias XbG_H630 : voltage is Vneg_temp(630);
	alias XbG_H631 : voltage is Vneg_temp(631);
	alias XbG_H632 : voltage is Vneg_temp(632);
	alias XbG_H633 : voltage is Vneg_temp(633);
	alias XbG_H634 : voltage is Vneg_temp(634);
	alias XbG_H635 : voltage is Vneg_temp(635);
	alias XbG_H636 : voltage is Vneg_temp(636);
	alias XbG_H637 : voltage is Vneg_temp(637);
	alias XbG_H638 : voltage is Vneg_temp(638);
	alias XbG_H639 : voltage is Vneg_temp(639);
	alias XbG_H640 : voltage is Vneg_temp(640);
	alias XbG_H641 : voltage is Vneg_temp(641);
	alias XbG_H642 : voltage is Vneg_temp(642);
	alias XbG_H643 : voltage is Vneg_temp(643);
	alias XbG_H644 : voltage is Vneg_temp(644);
	alias XbG_H645 : voltage is Vneg_temp(645);
	alias XbG_H646 : voltage is Vneg_temp(646);
	alias XbG_H647 : voltage is Vneg_temp(647);
	alias XbG_H648 : voltage is Vneg_temp(648);
	alias XbG_H649 : voltage is Vneg_temp(649);
	alias XbG_H650 : voltage is Vneg_temp(650);
	alias XbG_H651 : voltage is Vneg_temp(651);
	alias XbG_H652 : voltage is Vneg_temp(652);
	alias XbG_H653 : voltage is Vneg_temp(653);
	alias XbG_H654 : voltage is Vneg_temp(654);
	alias XbG_H655 : voltage is Vneg_temp(655);
	alias XbG_H656 : voltage is Vneg_temp(656);
	alias XbG_H657 : voltage is Vneg_temp(657);
	alias XbG_H658 : voltage is Vneg_temp(658);
	alias XbG_H659 : voltage is Vneg_temp(659);
	alias XbG_H660 : voltage is Vneg_temp(660);
	alias XbG_H661 : voltage is Vneg_temp(661);
	alias XbG_H662 : voltage is Vneg_temp(662);
	alias XbG_H663 : voltage is Vneg_temp(663);
	alias XbG_H664 : voltage is Vneg_temp(664);
	alias XbG_H665 : voltage is Vneg_temp(665);
	alias XbG_H666 : voltage is Vneg_temp(666);
	alias XbG_H667 : voltage is Vneg_temp(667);
	alias XbG_H668 : voltage is Vneg_temp(668);
	alias XbG_H669 : voltage is Vneg_temp(669);
	alias XbG_H670 : voltage is Vneg_temp(670);
	alias XbG_H671 : voltage is Vneg_temp(671);
	alias XbG_H672 : voltage is Vneg_temp(672);
	alias XbG_H673 : voltage is Vneg_temp(673);
	alias XbG_H674 : voltage is Vneg_temp(674);
	alias XbG_H675 : voltage is Vneg_temp(675);
	alias XbG_H676 : voltage is Vneg_temp(676);
	alias XbG_H677 : voltage is Vneg_temp(677);
	alias XbG_H678 : voltage is Vneg_temp(678);
	alias XbG_H679 : voltage is Vneg_temp(679);
	alias XbG_H680 : voltage is Vneg_temp(680);
	alias XbG_H681 : voltage is Vneg_temp(681);
	alias XbG_H682 : voltage is Vneg_temp(682);
	alias XbG_H683 : voltage is Vneg_temp(683);
	alias XbG_H684 : voltage is Vneg_temp(684);
	alias XbG_H685 : voltage is Vneg_temp(685);
	alias XbG_H686 : voltage is Vneg_temp(686);
	alias XbG_H687 : voltage is Vneg_temp(687);
	alias XbG_H688 : voltage is Vneg_temp(688);
	alias XbG_H689 : voltage is Vneg_temp(689);
	alias XbG_H690 : voltage is Vneg_temp(690);
	alias XbG_H691 : voltage is Vneg_temp(691);
	alias XbG_H692 : voltage is Vneg_temp(692);
	alias XbG_H693 : voltage is Vneg_temp(693);
	alias XbG_H694 : voltage is Vneg_temp(694);
	alias XbG_H695 : voltage is Vneg_temp(695);
	alias XbG_H696 : voltage is Vneg_temp(696);
	alias XbG_H697 : voltage is Vneg_temp(697);
	alias XbG_H698 : voltage is Vneg_temp(698);
	alias XbG_H699 : voltage is Vneg_temp(699);
	alias XbG_H700 : voltage is Vneg_temp(700);
	alias XbG_H701 : voltage is Vneg_temp(701);
	alias XbG_H702 : voltage is Vneg_temp(702);
	alias XbG_H703 : voltage is Vneg_temp(703);
	alias XbG_H704 : voltage is Vneg_temp(704);
	alias XbG_H705 : voltage is Vneg_temp(705);
	alias XbG_H706 : voltage is Vneg_temp(706);
	alias XbG_H707 : voltage is Vneg_temp(707);
	alias XbG_H708 : voltage is Vneg_temp(708);
	alias XbG_H709 : voltage is Vneg_temp(709);
	alias XbG_H710 : voltage is Vneg_temp(710);
	alias XbG_H711 : voltage is Vneg_temp(711);
	alias XbG_H712 : voltage is Vneg_temp(712);
	alias XbG_H713 : voltage is Vneg_temp(713);
	alias XbG_H714 : voltage is Vneg_temp(714);
	alias XbG_H715 : voltage is Vneg_temp(715);
	alias XbG_H716 : voltage is Vneg_temp(716);
	alias XbG_H717 : voltage is Vneg_temp(717);
	alias XbG_H718 : voltage is Vneg_temp(718);
	alias XbG_H719 : voltage is Vneg_temp(719);
	alias XbG_H720 : voltage is Vneg_temp(720);
	alias XbG_H721 : voltage is Vneg_temp(721);
	alias XbG_H722 : voltage is Vneg_temp(722);
	alias XbG_H723 : voltage is Vneg_temp(723);
	alias XbG_H724 : voltage is Vneg_temp(724);
	alias XbG_H725 : voltage is Vneg_temp(725);
	alias XbG_H726 : voltage is Vneg_temp(726);
	alias XbG_H727 : voltage is Vneg_temp(727);
	alias XbG_H728 : voltage is Vneg_temp(728);
	alias XbG_H729 : voltage is Vneg_temp(729);
	alias XbG_H730 : voltage is Vneg_temp(730);
	alias XbG_H731 : voltage is Vneg_temp(731);
	alias XbG_H732 : voltage is Vneg_temp(732);
	alias XbG_H733 : voltage is Vneg_temp(733);
	alias XbG_H734 : voltage is Vneg_temp(734);
	alias XbG_H735 : voltage is Vneg_temp(735);
alias po00_tmp : std_logic is output_temp(0);
alias po01_tmp : std_logic is output_temp(1);
alias po02_tmp : std_logic is output_temp(2);
alias po03_tmp : std_logic is output_temp(3);
alias po04_tmp : std_logic is output_temp(4);
alias po05_tmp : std_logic is output_temp(5);
alias po06_tmp : std_logic is output_temp(6);
alias po07_tmp : std_logic is output_temp(7);
alias po08_tmp : std_logic is output_temp(8);
alias po09_tmp : std_logic is output_temp(9);
alias po10_tmp : std_logic is output_temp(10);
alias po11_tmp : std_logic is output_temp(11);
alias po12_tmp : std_logic is output_temp(12);
alias po13_tmp : std_logic is output_temp(13);
alias po15_tmp : std_logic is output_temp(14);
alias po16_tmp : std_logic is output_temp(15);
alias po17_tmp : std_logic is output_temp(16);
alias po18_tmp : std_logic is output_temp(17);
alias po20_tmp : std_logic is output_temp(18);
alias po21_tmp : std_logic is output_temp(19);
alias po22_tmp : std_logic is output_temp(20);
alias po23_tmp : std_logic is output_temp(21);
alias po24_tmp : std_logic is output_temp(22);
alias po25_tmp : std_logic is output_temp(23);
alias po26_tmp : std_logic is output_temp(24);
alias po27_tmp : std_logic is output_temp(25);
alias po28_tmp : std_logic is output_temp(26);
alias po29_tmp : std_logic is output_temp(27);
alias po30_tmp : std_logic is output_temp(28);
alias po31_tmp : std_logic is output_temp(29);
alias po32_tmp : std_logic is output_temp(30);
alias po33_tmp : std_logic is output_temp(31);
alias po34_tmp : std_logic is output_temp(32);
alias po35_tmp : std_logic is output_temp(33);
alias po36_tmp : std_logic is output_temp(34);
alias po37_tmp : std_logic is output_temp(35);
alias po38_tmp : std_logic is output_temp(36);
alias po39_tmp : std_logic is output_temp(37);
alias po40_tmp : std_logic is output_temp(38);
alias po41_tmp : std_logic is output_temp(39);
alias po42_tmp : std_logic is output_temp(40);
alias po43_tmp : std_logic is output_temp(41);
alias po44_tmp : std_logic is output_temp(42);
alias po45_tmp : std_logic is output_temp(43);
alias po46_tmp : std_logic is output_temp(44);
alias po47_tmp : std_logic is output_temp(45);
alias po48_tmp : std_logic is output_temp(46);
alias po49_tmp : std_logic is output_temp(47);
alias po50_tmp : std_logic is output_temp(48);
alias po51_tmp : std_logic is output_temp(49);
alias po52_tmp : std_logic is output_temp(50);
alias po53_tmp : std_logic is output_temp(51);
alias po54_tmp : std_logic is output_temp(52);
alias po55_tmp : std_logic is output_temp(53);
alias li0_tmp : std_logic is output_temp(54);
alias li1_tmp : std_logic is output_temp(55);
alias li2_tmp : std_logic is output_temp(56);
alias li3_tmp : std_logic is output_temp(57);
alias li4_tmp : std_logic is output_temp(58);
alias li5_tmp : std_logic is output_temp(59);
alias li6_tmp : std_logic is output_temp(60);
type FSMstate is (IDLE,A_INA,B_RI,C_CFM,D_EVM,E_EVR,F_INR,G_SS);

signal state, next_state : FSMstate := IDLE;

signal feedback_enable : std_logic := '0';
signal current_state: std_logic_vector(6 downto 0) := (others=>'0');
signal clk : std_logic := '0';

constant clk_period : time := 1 ns;

function vectorize(V: std_logic) return std_logic_vector is
variable v_tmp : std_logic_vector(0 downto 0);
begin
v_tmp(0) := V;
return v_tmp;
end vectorize;

begin

Inst_Crossbar : crossbar_1 PORT MAP(
Vpos => Vpos_temp,
Vneg => Vneg_temp,
output => output_temp
);

po00<=po00_tmp;
po01<=po01_tmp;
po02<=po02_tmp;
po03<=po03_tmp;
po04<=po04_tmp;
po05<=po05_tmp;
po06<=po06_tmp;
po07<=po07_tmp;
po08<=po08_tmp;
po09<=po09_tmp;
po10<=po10_tmp;
po11<=po11_tmp;
po12<=po12_tmp;
po13<=po13_tmp;
po15<=po15_tmp;
po16<=po16_tmp;
po17<=po17_tmp;
po18<=po18_tmp;
po20<=po20_tmp;
po21<=po21_tmp;
po22<=po22_tmp;
po23<=po23_tmp;
po24<=po24_tmp;
po25<=po25_tmp;
po26<=po26_tmp;
po27<=po27_tmp;
po28<=po28_tmp;
po29<=po29_tmp;
po30<=po30_tmp;
po31<=po31_tmp;
po32<=po32_tmp;
po33<=po33_tmp;
po34<=po34_tmp;
po35<=po35_tmp;
po36<=po36_tmp;
po37<=po37_tmp;
po38<=po38_tmp;
po39<=po39_tmp;
po40<=po40_tmp;
po41<=po41_tmp;
po42<=po42_tmp;
po43<=po43_tmp;
po44<=po44_tmp;
po45<=po45_tmp;
po46<=po46_tmp;
po47<=po47_tmp;
po48<=po48_tmp;
po49<=po49_tmp;
po50<=po50_tmp;
po51<=po51_tmp;
po52<=po52_tmp;
po53<=po53_tmp;
po54<=po54_tmp;
po55<=po55_tmp;
li0<=li0_tmp;
li1<=li1_tmp;
li2<=li2_tmp;
li3<=li3_tmp;
li4<=li4_tmp;
li5<=li5_tmp;
li6<=li6_tmp;

-- Clock process definitions
clk_process : process (clk)
begin
clk <= not(clk) after clk_period/2; --only behavioral simulation
end process;

change_state: process (clk)
begin
if(clk'event and clk='1') then
state <= next_state;   --state change.
end if;
end process;

FSM: process(state,pi26,pi15,lo6,lo5,lo4,lo3,lo2,lo1,lo0,pi00,pi06,pi03,pi07,pi08,pi09,pi10,pi02,pi17,pi01,pi11,pi12,pi13,pi14,pi04,pi16,pi05,pi18,pi19,pi20,pi21,pi22,pi23,pi24,pi25,en)
begin

case state is

when IDLE =>

XbG_H0<=Vr;
XbG_H1<=Vr;
XbG_H10<=Vr;
XbG_H100<=Vr;
XbG_H101<=Vr;
XbG_H102<=Vr;
XbG_H103<=Vr;
XbG_H104<=Vr;
XbG_H105<=Vr;
XbG_H106<=Vr;
XbG_H107<=Vr;
XbG_H108<=Vr;
XbG_H109<=Vr;
XbG_H11<=Vr;
XbG_H110<=Vr;
XbG_H111<=Vr;
XbG_H112<=Vr;
XbG_H113<=Vr;
XbG_H114<=Vr;
XbG_H115<=Vr;
XbG_H116<=Vr;
XbG_H117<=Vr;
XbG_H118<=Vr;
XbG_H119<=Vr;
XbG_H12<=Vr;
XbG_H120<=Vr;
XbG_H121<=Vr;
XbG_H122<=Vr;
XbG_H123<=Vr;
XbG_H124<=Vr;
XbG_H125<=Vr;
XbG_H126<=Vr;
XbG_H127<=Vr;
XbG_H128<=Vr;
XbG_H129<=Vr;
XbG_H13<=Vr;
XbG_H130<=Vr;
XbG_H131<=Vr;
XbG_H132<=Vr;
XbG_H133<=Vr;
XbG_H134<=Vr;
XbG_H135<=Vr;
XbG_H136<=Vr;
XbG_H137<=Vr;
XbG_H138<=Vr;
XbG_H139<=Vr;
XbG_H14<=Vr;
XbG_H140<=Vr;
XbG_H141<=Vr;
XbG_H142<=Vr;
XbG_H143<=Vr;
XbG_H144<=Vr;
XbG_H145<=Vr;
XbG_H146<=Vr;
XbG_H147<=Vr;
XbG_H148<=Vr;
XbG_H149<=Vr;
XbG_H15<=Vr;
XbG_H150<=Vr;
XbG_H151<=Vr;
XbG_H152<=Vr;
XbG_H153<=Vr;
XbG_H154<=Vr;
XbG_H155<=Vr;
XbG_H156<=Vr;
XbG_H157<=Vr;
XbG_H158<=Vr;
XbG_H159<=Vr;
XbG_H16<=Vr;
XbG_H160<=Vr;
XbG_H161<=Vr;
XbG_H162<=Vr;
XbG_H163<=Vr;
XbG_H164<=Vr;
XbG_H165<=Vr;
XbG_H166<=Vr;
XbG_H167<=Vr;
XbG_H168<=Vr;
XbG_H169<=Vr;
XbG_H17<=Vr;
XbG_H170<=Vr;
XbG_H171<=Vr;
XbG_H172<=Vr;
XbG_H173<=Vr;
XbG_H174<=Vr;
XbG_H175<=Vr;
XbG_H176<=Vr;
XbG_H177<=Vr;
XbG_H178<=Vr;
XbG_H179<=Vr;
XbG_H18<=Vr;
XbG_H180<=Vr;
XbG_H181<=Vr;
XbG_H182<=Vr;
XbG_H183<=Vr;
XbG_H184<=Vr;
XbG_H185<=Vr;
XbG_H186<=Vr;
XbG_H187<=Vr;
XbG_H188<=Vr;
XbG_H189<=Vr;
XbG_H19<=Vr;
XbG_H190<=Vr;
XbG_H191<=Vr;
XbG_H192<=Vr;
XbG_H193<=Vr;
XbG_H194<=Vr;
XbG_H195<=Vr;
XbG_H196<=Vr;
XbG_H197<=Vr;
XbG_H198<=Vr;
XbG_H199<=Vr;
XbG_H2<=Vr;
XbG_H20<=Vr;
XbG_H200<=Vr;
XbG_H201<=Vr;
XbG_H202<=Vr;
XbG_H203<=Vr;
XbG_H204<=Vr;
XbG_H205<=Vr;
XbG_H206<=Vr;
XbG_H207<=Vr;
XbG_H208<=Vr;
XbG_H209<=Vr;
XbG_H21<=Vr;
XbG_H210<=Vr;
XbG_H211<=Vr;
XbG_H212<=Vr;
XbG_H213<=Vr;
XbG_H214<=Vr;
XbG_H215<=Vr;
XbG_H216<=Vr;
XbG_H217<=Vr;
XbG_H218<=Vr;
XbG_H219<=Vr;
XbG_H22<=Vr;
XbG_H220<=Vr;
XbG_H221<=Vr;
XbG_H222<=Vr;
XbG_H223<=Vr;
XbG_H224<=Vr;
XbG_H225<=Vr;
XbG_H226<=Vr;
XbG_H227<=Vr;
XbG_H228<=Vr;
XbG_H229<=Vr;
XbG_H23<=Vr;
XbG_H230<=Vr;
XbG_H231<=Vr;
XbG_H232<=Vr;
XbG_H233<=Vr;
XbG_H234<=Vr;
XbG_H235<=Vr;
XbG_H236<=Vr;
XbG_H237<=Vr;
XbG_H238<=Vr;
XbG_H239<=Vr;
XbG_H24<=Vr;
XbG_H240<=Vr;
XbG_H241<=Vr;
XbG_H242<=Vr;
XbG_H243<=Vr;
XbG_H244<=Vr;
XbG_H245<=Vr;
XbG_H246<=Vr;
XbG_H247<=Vr;
XbG_H248<=Vr;
XbG_H249<=Vr;
XbG_H25<=Vr;
XbG_H250<=Vr;
XbG_H251<=Vr;
XbG_H252<=Vr;
XbG_H253<=Vr;
XbG_H254<=Vr;
XbG_H255<=Vr;
XbG_H256<=Vr;
XbG_H257<=Vr;
XbG_H258<=Vr;
XbG_H259<=Vr;
XbG_H26<=Vr;
XbG_H260<=Vr;
XbG_H261<=Vr;
XbG_H262<=Vr;
XbG_H263<=Vr;
XbG_H264<=Vr;
XbG_H265<=Vr;
XbG_H266<=Vr;
XbG_H267<=Vr;
XbG_H268<=Vr;
XbG_H269<=Vr;
XbG_H27<=Vr;
XbG_H270<=Vr;
XbG_H271<=Vr;
XbG_H272<=Vr;
XbG_H273<=Vr;
XbG_H274<=Vr;
XbG_H275<=Vr;
XbG_H276<=Vr;
XbG_H277<=Vr;
XbG_H278<=Vr;
XbG_H279<=Vr;
XbG_H28<=Vr;
XbG_H280<=Vr;
XbG_H281<=Vr;
XbG_H282<=Vr;
XbG_H283<=Vr;
XbG_H284<=Vr;
XbG_H285<=Vr;
XbG_H286<=Vr;
XbG_H287<=Vr;
XbG_H288<=Vr;
XbG_H289<=Vr;
XbG_H29<=Vr;
XbG_H290<=Vr;
XbG_H291<=Vr;
XbG_H292<=Vr;
XbG_H293<=Vr;
XbG_H294<=Vr;
XbG_H295<=Vr;
XbG_H296<=Vr;
XbG_H297<=Vr;
XbG_H298<=Vr;
XbG_H299<=Vr;
XbG_H3<=Vr;
XbG_H30<=Vr;
XbG_H300<=Vr;
XbG_H301<=Vr;
XbG_H302<=Vr;
XbG_H303<=Vr;
XbG_H304<=Vr;
XbG_H305<=Vr;
XbG_H306<=Vr;
XbG_H307<=Vr;
XbG_H308<=Vr;
XbG_H309<=Vr;
XbG_H31<=Vr;
XbG_H310<=Vr;
XbG_H311<=Vr;
XbG_H312<=Vr;
XbG_H313<=Vr;
XbG_H314<=Vr;
XbG_H315<=Vr;
XbG_H316<=Vr;
XbG_H317<=Vr;
XbG_H318<=Vr;
XbG_H319<=Vr;
XbG_H32<=Vr;
XbG_H320<=Vr;
XbG_H321<=Vr;
XbG_H322<=Vr;
XbG_H323<=Vr;
XbG_H324<=Vr;
XbG_H325<=Vr;
XbG_H326<=Vr;
XbG_H327<=Vr;
XbG_H328<=Vr;
XbG_H329<=Vr;
XbG_H33<=Vr;
XbG_H330<=Vr;
XbG_H331<=Vr;
XbG_H332<=Vr;
XbG_H333<=Vr;
XbG_H334<=Vr;
XbG_H335<=Vr;
XbG_H336<=Vr;
XbG_H337<=Vr;
XbG_H338<=Vr;
XbG_H339<=Vr;
XbG_H34<=Vr;
XbG_H340<=Vr;
XbG_H341<=Vr;
XbG_H342<=Vr;
XbG_H343<=Vr;
XbG_H344<=Vr;
XbG_H345<=Vr;
XbG_H346<=Vr;
XbG_H347<=Vr;
XbG_H348<=Vr;
XbG_H349<=Vr;
XbG_H35<=Vr;
XbG_H350<=Vr;
XbG_H351<=Vr;
XbG_H352<=Vr;
XbG_H353<=Vr;
XbG_H354<=Vr;
XbG_H355<=Vr;
XbG_H356<=Vr;
XbG_H357<=Vr;
XbG_H358<=Vr;
XbG_H359<=Vr;
XbG_H36<=Vr;
XbG_H360<=Vr;
XbG_H361<=Vr;
XbG_H362<=Vr;
XbG_H363<=Vr;
XbG_H364<=Vr;
XbG_H365<=Vr;
XbG_H366<=Vr;
XbG_H367<=Vr;
XbG_H368<=Vr;
XbG_H369<=Vr;
XbG_H37<=Vr;
XbG_H370<=Vr;
XbG_H371<=Vr;
XbG_H372<=Vr;
XbG_H373<=Vr;
XbG_H374<=Vr;
XbG_H375<=Vr;
XbG_H376<=Vr;
XbG_H377<=Vr;
XbG_H378<=Vr;
XbG_H379<=Vr;
XbG_H38<=Vr;
XbG_H380<=Vr;
XbG_H381<=Vr;
XbG_H382<=Vr;
XbG_H383<=Vr;
XbG_H384<=Vr;
XbG_H385<=Vr;
XbG_H386<=Vr;
XbG_H387<=Vr;
XbG_H388<=Vr;
XbG_H389<=Vr;
XbG_H39<=Vr;
XbG_H390<=Vr;
XbG_H391<=Vr;
XbG_H392<=Vr;
XbG_H393<=Vr;
XbG_H394<=Vr;
XbG_H395<=Vr;
XbG_H396<=Vr;
XbG_H397<=Vr;
XbG_H398<=Vr;
XbG_H399<=Vr;
XbG_H4<=Vr;
XbG_H40<=Vr;
XbG_H400<=Vr;
XbG_H401<=Vr;
XbG_H402<=Vr;
XbG_H403<=Vr;
XbG_H404<=Vr;
XbG_H405<=Vr;
XbG_H406<=Vr;
XbG_H407<=Vr;
XbG_H408<=Vr;
XbG_H409<=Vr;
XbG_H41<=Vr;
XbG_H410<=Vr;
XbG_H411<=Vr;
XbG_H412<=Vr;
XbG_H413<=Vr;
XbG_H414<=Vr;
XbG_H415<=Vr;
XbG_H416<=Vr;
XbG_H417<=Vr;
XbG_H418<=Vr;
XbG_H419<=Vr;
XbG_H42<=Vr;
XbG_H420<=Vr;
XbG_H421<=Vr;
XbG_H422<=Vr;
XbG_H423<=Vr;
XbG_H424<=Vr;
XbG_H425<=Vr;
XbG_H426<=Vr;
XbG_H427<=Vr;
XbG_H428<=Vr;
XbG_H429<=Vr;
XbG_H43<=Vr;
XbG_H430<=Vr;
XbG_H431<=Vr;
XbG_H432<=Vr;
XbG_H433<=Vr;
XbG_H434<=Vr;
XbG_H435<=Vr;
XbG_H436<=Vr;
XbG_H437<=Vr;
XbG_H438<=Vr;
XbG_H439<=Vr;
XbG_H44<=Vr;
XbG_H440<=Vr;
XbG_H441<=Vr;
XbG_H442<=Vr;
XbG_H443<=Vr;
XbG_H444<=Vr;
XbG_H445<=Vr;
XbG_H446<=Vr;
XbG_H447<=Vr;
XbG_H448<=Vr;
XbG_H449<=Vr;
XbG_H45<=Vr;
XbG_H450<=Vr;
XbG_H451<=Vr;
XbG_H452<=Vr;
XbG_H453<=Vr;
XbG_H454<=Vr;
XbG_H455<=Vr;
XbG_H456<=Vr;
XbG_H457<=Vr;
XbG_H458<=Vr;
XbG_H459<=Vr;
XbG_H46<=Vr;
XbG_H460<=Vr;
XbG_H461<=Vr;
XbG_H462<=Vr;
XbG_H463<=Vr;
XbG_H464<=Vr;
XbG_H465<=Vr;
XbG_H466<=Vr;
XbG_H467<=Vr;
XbG_H468<=Vr;
XbG_H469<=Vr;
XbG_H47<=Vr;
XbG_H470<=Vr;
XbG_H471<=Vr;
XbG_H472<=Vr;
XbG_H473<=Vr;
XbG_H474<=Vr;
XbG_H475<=Vr;
XbG_H476<=Vr;
XbG_H477<=Vr;
XbG_H478<=Vr;
XbG_H479<=Vr;
XbG_H48<=Vr;
XbG_H480<=Vr;
XbG_H481<=Vr;
XbG_H482<=Vr;
XbG_H483<=Vr;
XbG_H484<=Vr;
XbG_H485<=Vr;
XbG_H486<=Vr;
XbG_H487<=Vr;
XbG_H488<=Vr;
XbG_H489<=Vr;
XbG_H49<=Vr;
XbG_H490<=Vr;
XbG_H491<=Vr;
XbG_H492<=Vr;
XbG_H493<=Vr;
XbG_H494<=Vr;
XbG_H495<=Vr;
XbG_H496<=Vr;
XbG_H497<=Vr;
XbG_H498<=Vr;
XbG_H499<=Vr;
XbG_H5<=Vr;
XbG_H50<=Vr;
XbG_H500<=Vr;
XbG_H501<=Vr;
XbG_H502<=Vr;
XbG_H503<=Vr;
XbG_H504<=Vr;
XbG_H505<=Vr;
XbG_H506<=Vr;
XbG_H507<=Vr;
XbG_H508<=Vr;
XbG_H509<=Vr;
XbG_H51<=Vr;
XbG_H510<=Vr;
XbG_H511<=Vr;
XbG_H512<=Vr;
XbG_H513<=Vr;
XbG_H514<=Vr;
XbG_H515<=Vr;
XbG_H516<=Vr;
XbG_H517<=Vr;
XbG_H518<=Vr;
XbG_H519<=Vr;
XbG_H52<=Vr;
XbG_H520<=Vr;
XbG_H521<=Vr;
XbG_H522<=Vr;
XbG_H523<=Vr;
XbG_H524<=Vr;
XbG_H525<=Vr;
XbG_H526<=Vr;
XbG_H527<=Vr;
XbG_H528<=Vr;
XbG_H529<=Vr;
XbG_H53<=Vr;
XbG_H530<=Vr;
XbG_H531<=Vr;
XbG_H532<=Vr;
XbG_H533<=Vr;
XbG_H534<=Vr;
XbG_H535<=Vr;
XbG_H536<=Vr;
XbG_H537<=Vr;
XbG_H538<=Vr;
XbG_H539<=Vr;
XbG_H54<=Vr;
XbG_H540<=Vr;
XbG_H541<=Vr;
XbG_H542<=Vr;
XbG_H543<=Vr;
XbG_H544<=Vr;
XbG_H545<=Vr;
XbG_H546<=Vr;
XbG_H547<=Vr;
XbG_H548<=Vr;
XbG_H549<=Vr;
XbG_H55<=Vr;
XbG_H550<=Vr;
XbG_H551<=Vr;
XbG_H552<=Vr;
XbG_H553<=Vr;
XbG_H554<=Vr;
XbG_H555<=Vr;
XbG_H556<=Vr;
XbG_H557<=Vr;
XbG_H558<=Vr;
XbG_H559<=Vr;
XbG_H56<=Vr;
XbG_H560<=Vr;
XbG_H561<=Vr;
XbG_H562<=Vr;
XbG_H563<=Vr;
XbG_H564<=Vr;
XbG_H565<=Vr;
XbG_H566<=Vr;
XbG_H567<=Vr;
XbG_H568<=Vr;
XbG_H569<=Vr;
XbG_H57<=Vr;
XbG_H570<=Vr;
XbG_H571<=Vr;
XbG_H572<=Vr;
XbG_H573<=Vr;
XbG_H574<=Vr;
XbG_H575<=Vr;
XbG_H576<=Vr;
XbG_H577<=Vr;
XbG_H578<=Vr;
XbG_H579<=Vr;
XbG_H58<=Vr;
XbG_H580<=Vr;
XbG_H581<=Vr;
XbG_H582<=Vr;
XbG_H583<=Vr;
XbG_H584<=Vr;
XbG_H585<=Vr;
XbG_H586<=Vr;
XbG_H587<=Vr;
XbG_H588<=Vr;
XbG_H589<=Vr;
XbG_H59<=Vr;
XbG_H590<=Vr;
XbG_H591<=Vr;
XbG_H592<=Vr;
XbG_H593<=Vr;
XbG_H594<=Vr;
XbG_H595<=Vr;
XbG_H596<=Vr;
XbG_H597<=Vr;
XbG_H598<=Vr;
XbG_H599<=Vr;
XbG_H6<=Vr;
XbG_H60<=Vr;
XbG_H600<=Vr;
XbG_H601<=Vr;
XbG_H602<=Vr;
XbG_H603<=Vr;
XbG_H604<=Vr;
XbG_H605<=Vr;
XbG_H606<=Vr;
XbG_H607<=Vr;
XbG_H608<=Vr;
XbG_H609<=Vr;
XbG_H61<=Vr;
XbG_H610<=Vr;
XbG_H611<=Vr;
XbG_H612<=Vr;
XbG_H613<=Vr;
XbG_H614<=Vr;
XbG_H615<=Vr;
XbG_H616<=Vr;
XbG_H617<=Vr;
XbG_H618<=Vr;
XbG_H619<=Vr;
XbG_H62<=Vr;
XbG_H620<=Vr;
XbG_H621<=Vr;
XbG_H622<=Vr;
XbG_H623<=Vr;
XbG_H624<=Vr;
XbG_H625<=Vr;
XbG_H626<=Vr;
XbG_H627<=Vr;
XbG_H628<=Vr;
XbG_H629<=Vr;
XbG_H63<=Vr;
XbG_H630<=Vr;
XbG_H631<=Vr;
XbG_H632<=Vr;
XbG_H633<=Vr;
XbG_H634<=Vr;
XbG_H635<=Vr;
XbG_H636<=Vr;
XbG_H637<=Vr;
XbG_H638<=Vr;
XbG_H639<=Vr;
XbG_H64<=Vr;
XbG_H640<=Vr;
XbG_H641<=Vr;
XbG_H642<=Vr;
XbG_H643<=Vr;
XbG_H644<=Vr;
XbG_H645<=Vr;
XbG_H646<=Vr;
XbG_H647<=Vr;
XbG_H648<=Vr;
XbG_H649<=Vr;
XbG_H65<=Vr;
XbG_H650<=Vr;
XbG_H651<=Vr;
XbG_H652<=Vr;
XbG_H653<=Vr;
XbG_H654<=Vr;
XbG_H655<=Vr;
XbG_H656<=Vr;
XbG_H657<=Vr;
XbG_H658<=Vr;
XbG_H659<=Vr;
XbG_H66<=Vr;
XbG_H660<=Vr;
XbG_H661<=Vr;
XbG_H662<=Vr;
XbG_H663<=Vr;
XbG_H664<=Vr;
XbG_H665<=Vr;
XbG_H666<=Vr;
XbG_H667<=Vr;
XbG_H668<=Vr;
XbG_H669<=Vr;
XbG_H67<=Vr;
XbG_H670<=Vr;
XbG_H671<=Vr;
XbG_H672<=Vr;
XbG_H673<=Vr;
XbG_H674<=Vr;
XbG_H675<=Vr;
XbG_H676<=Vr;
XbG_H677<=Vr;
XbG_H678<=Vr;
XbG_H679<=Vr;
XbG_H68<=Vr;
XbG_H680<=Vr;
XbG_H681<=Vr;
XbG_H682<=Vr;
XbG_H683<=Vr;
XbG_H684<=Vr;
XbG_H685<=Vr;
XbG_H686<=Vr;
XbG_H687<=Vr;
XbG_H688<=Vr;
XbG_H689<=Vr;
XbG_H69<=Vr;
XbG_H690<=Vr;
XbG_H691<=Vr;
XbG_H692<=Vr;
XbG_H693<=Vr;
XbG_H694<=Vr;
XbG_H695<=Vr;
XbG_H696<=Vr;
XbG_H697<=Vr;
XbG_H698<=Vr;
XbG_H699<=Vr;
XbG_H7<=Vr;
XbG_H70<=Vr;
XbG_H700<=Vr;
XbG_H701<=Vr;
XbG_H702<=Vr;
XbG_H703<=Vr;
XbG_H704<=Vr;
XbG_H705<=Vr;
XbG_H706<=Vr;
XbG_H707<=Vr;
XbG_H708<=Vr;
XbG_H709<=Vr;
XbG_H71<=Vr;
XbG_H710<=Vr;
XbG_H711<=Vr;
XbG_H712<=Vr;
XbG_H713<=Vr;
XbG_H714<=Vr;
XbG_H715<=Vr;
XbG_H716<=Vr;
XbG_H717<=Vr;
XbG_H718<=Vr;
XbG_H719<=Vr;
XbG_H72<=Vr;
XbG_H720<=Vr;
XbG_H721<=Vr;
XbG_H722<=Vr;
XbG_H723<=Vr;
XbG_H724<=Vr;
XbG_H725<=Vr;
XbG_H726<=Vr;
XbG_H727<=Vr;
XbG_H728<=Vr;
XbG_H729<=Vr;
XbG_H73<=Vr;
XbG_H730<=Vr;
XbG_H731<=Vr;
XbG_H732<=Vr;
XbG_H733<=Vr;
XbG_H734<=Vr;
XbG_H735<=Vr;
XbG_H74<=Vr;
XbG_H75<=Vr;
XbG_H76<=Vr;
XbG_H77<=Vr;
XbG_H78<=Vr;
XbG_H79<=Vr;
XbG_H8<=Vr;
XbG_H80<=Vr;
XbG_H81<=Vr;
XbG_H82<=Vr;
XbG_H83<=Vr;
XbG_H84<=Vr;
XbG_H85<=Vr;
XbG_H86<=Vr;
XbG_H87<=Vr;
XbG_H88<=Vr;
XbG_H89<=Vr;
XbG_H9<=Vr;
XbG_H90<=Vr;
XbG_H91<=Vr;
XbG_H92<=Vr;
XbG_H93<=Vr;
XbG_H94<=Vr;
XbG_H95<=Vr;
XbG_H96<=Vr;
XbG_H97<=Vr;
XbG_H98<=Vr;
XbG_H99<=Vr;
XbG_V0<=Vr;
XbG_V1<=Vr;
XbG_V10<=Vr;
XbG_V100<=Vr;
XbG_V101<=Vr;
XbG_V102<=Vr;
XbG_V103<=Vr;
XbG_V104<=Vr;
XbG_V105<=Vr;
XbG_V106<=Vr;
XbG_V107<=Vr;
XbG_V108<=Vr;
XbG_V109<=Vr;
XbG_V11<=Vr;
XbG_V110<=Vr;
XbG_V111<=Vr;
XbG_V112<=Vr;
XbG_V113<=Vr;
XbG_V114<=Vr;
XbG_V115<=Vr;
XbG_V116<=Vr;
XbG_V117<=Vr;
XbG_V118<=Vr;
XbG_V119<=Vr;
XbG_V12<=Vr;
XbG_V120<=Vr;
XbG_V121<=Vr;
XbG_V122<=Vr;
XbG_V123<=Vr;
XbG_V124<=Vr;
XbG_V125<=Vr;
XbG_V126<=Vr;
XbG_V127<=Vr;
XbG_V128<=Vr;
XbG_V129<=Vr;
XbG_V13<=Vr;
XbG_V130<=Vr;
XbG_V131<=Vr;
XbG_V132<=Vr;
XbG_V133<=Vr;
XbG_V134<=Vr;
XbG_V135<=Vr;
XbG_V136<=Vr;
XbG_V137<=Vr;
XbG_V138<=Vr;
XbG_V139<=Vr;
XbG_V14<=Vr;
XbG_V140<=Vr;
XbG_V141<=Vr;
XbG_V142<=Vr;
XbG_V143<=Vr;
XbG_V144<=Vr;
XbG_V145<=Vr;
XbG_V146<=Vr;
XbG_V147<=Vr;
XbG_V148<=Vr;
XbG_V149<=Vr;
XbG_V15<=Vr;
XbG_V150<=Vr;
XbG_V151<=Vr;
XbG_V152<=Vr;
XbG_V153<=Vr;
XbG_V154<=Vr;
XbG_V155<=Vr;
XbG_V156<=Vr;
XbG_V157<=Vr;
XbG_V158<=Vr;
XbG_V159<=Vr;
XbG_V16<=Vr;
XbG_V160<=Vr;
XbG_V161<=Vr;
XbG_V162<=Vr;
XbG_V163<=Vr;
XbG_V164<=Vr;
XbG_V165<=Vr;
XbG_V166<=Vr;
XbG_V167<=Vr;
XbG_V168<=Vr;
XbG_V169<=Vr;
XbG_V17<=Vr;
XbG_V170<=Vr;
XbG_V171<=Vr;
XbG_V172<=Vr;
XbG_V173<=Vr;
XbG_V174<=Vr;
XbG_V175<=Vr;
XbG_V176<=Vr;
XbG_V177<=Vr;
XbG_V178<=Vr;
XbG_V179<=Vr;
XbG_V18<=Vr;
XbG_V180<=Vr;
XbG_V181<=Vr;
XbG_V182<=Vr;
XbG_V183<=Vr;
XbG_V184<=Vr;
XbG_V185<=Vr;
XbG_V186<=Vr;
XbG_V187<=Vr;
XbG_V188<=Vr;
XbG_V189<=Vr;
XbG_V19<=Vr;
XbG_V2<=Vr;
XbG_V20<=Vr;
XbG_V21<=Vr;
XbG_V22<=Vr;
XbG_V23<=Vr;
XbG_V24<=Vr;
XbG_V25<=Vr;
XbG_V26<=Vr;
XbG_V27<=Vr;
XbG_V28<=Vr;
XbG_V29<=Vr;
XbG_V3<=Vr;
XbG_V30<=Vr;
XbG_V31<=Vr;
XbG_V32<=Vr;
XbG_V33<=Vr;
XbG_V34<=Vr;
XbG_V35<=Vr;
XbG_V36<=Vr;
XbG_V37<=Vr;
XbG_V38<=Vr;
XbG_V39<=Vr;
XbG_V4<=Vr;
XbG_V40<=Vr;
XbG_V41<=Vr;
XbG_V42<=Vr;
XbG_V43<=Vr;
XbG_V44<=Vr;
XbG_V45<=Vr;
XbG_V46<=Vr;
XbG_V47<=Vr;
XbG_V48<=Vr;
XbG_V49<=Vr;
XbG_V5<=Vr;
XbG_V50<=Vr;
XbG_V51<=Vr;
XbG_V52<=Vr;
XbG_V53<=Vr;
XbG_V54<=Vr;
XbG_V55<=Vr;
XbG_V56<=Vr;
XbG_V57<=Vr;
XbG_V58<=Vr;
XbG_V59<=Vr;
XbG_V6<=Vr;
XbG_V60<=Vr;
XbG_V61<=Vr;
XbG_V62<=Vr;
XbG_V63<=Vr;
XbG_V64<=Vr;
XbG_V65<=Vr;
XbG_V66<=Vr;
XbG_V67<=Vr;
XbG_V68<=Vr;
XbG_V69<=Vr;
XbG_V7<=Vr;
XbG_V70<=Vr;
XbG_V71<=Vr;
XbG_V72<=Vr;
XbG_V73<=Vr;
XbG_V74<=Vr;
XbG_V75<=Vr;
XbG_V76<=Vr;
XbG_V77<=Vr;
XbG_V78<=Vr;
XbG_V79<=Vr;
XbG_V8<=Vr;
XbG_V80<=Vr;
XbG_V81<=Vr;
XbG_V82<=Vr;
XbG_V83<=Vr;
XbG_V84<=Vr;
XbG_V85<=Vr;
XbG_V86<=Vr;
XbG_V87<=Vr;
XbG_V88<=Vr;
XbG_V89<=Vr;
XbG_V9<=Vr;
XbG_V90<=Vr;
XbG_V91<=Vr;
XbG_V92<=Vr;
XbG_V93<=Vr;
XbG_V94<=Vr;
XbG_V95<=Vr;
XbG_V96<=Vr;
XbG_V97<=Vr;
XbG_V98<=Vr;
XbG_V99<=Vr;
if feedback_enable = '0' then
current_state(6 downto 0) <= vectorize(lo0)&vectorize(lo1)&vectorize(lo2)&vectorize(lo3)&vectorize(lo4)&vectorize(lo5)&vectorize(lo6);
else
current_state(6 downto 0) <= vectorize(li0_tmp)&vectorize(li1_tmp)&vectorize(li2_tmp)&vectorize(li3_tmp)&vectorize(li4_tmp)&vectorize(li5_tmp)&vectorize(li6_tmp);
end if;

done<='0' after clk_period;

if(en='1') then
next_state<=A_INA;
else
next_state<=IDLE;
end if;

when A_INA =>


if feedback_enable = '0' then

XbG_H0<=Vw;
XbG_H1<=Vw;
XbG_H10<=Vw;
XbG_H100<=Vw;
XbG_H101<=Vw;
XbG_H102<=Vw;
XbG_H103<=Vw;
XbG_H104<=Vw;
XbG_H105<=Vw;
XbG_H106<=Vw;
XbG_H107<=Vw;
XbG_H108<=Vw;
XbG_H109<=Vw;
XbG_H11<=Vw;
XbG_H110<=Vw;
XbG_H111<=Vw;
XbG_H112<=Vw;
XbG_H113<=Vw;
XbG_H114<=Vw;
XbG_H115<=Vw;
XbG_H116<=Vw;
XbG_H117<=Vw;
XbG_H118<=Vw;
XbG_H119<=Vw;
XbG_H12<=Vw;
XbG_H120<=Vw;
XbG_H121<=Vw;
XbG_H122<=Vw;
XbG_H123<=Vw;
XbG_H124<=Vw;
XbG_H125<=Vw;
XbG_H126<=Vw;
XbG_H127<=Vw;
XbG_H128<=Vw;
XbG_H129<=Vw;
XbG_H13<=Vw;
XbG_H130<=Vw;
XbG_H131<=Vw;
XbG_H132<=Vw;
XbG_H133<=Vw;
XbG_H134<=Vw;
XbG_H135<=Vw;
XbG_H136<=Vw;
XbG_H137<=Vw;
XbG_H138<=Vw;
XbG_H139<=Vw;
XbG_H14<=Vw;
XbG_H140<=Vw;
XbG_H141<=Vw;
XbG_H142<=Vw;
XbG_H143<=Vw;
XbG_H144<=Vw;
XbG_H145<=Vw;
XbG_H146<=Vw;
XbG_H147<=Vw;
XbG_H148<=Vw;
XbG_H149<=Vw;
XbG_H15<=Vw;
XbG_H150<=Vw;
XbG_H151<=Vw;
XbG_H152<=Vw;
XbG_H153<=Vw;
XbG_H154<=Vw;
XbG_H155<=Vw;
XbG_H156<=Vw;
XbG_H157<=Vw;
XbG_H158<=Vw;
XbG_H159<=Vw;
XbG_H16<=Vw;
XbG_H160<=Vw;
XbG_H161<=Vw;
XbG_H162<=Vw;
XbG_H163<=Vw;
XbG_H164<=Vw;
XbG_H165<=Vw;
XbG_H166<=Vw;
XbG_H167<=Vw;
XbG_H168<=Vw;
XbG_H169<=Vw;
XbG_H17<=Vw;
XbG_H170<=Vw;
XbG_H171<=Vw;
XbG_H172<=Vw;
XbG_H173<=Vw;
XbG_H174<=Vw;
XbG_H175<=Vw;
XbG_H176<=Vw;
XbG_H177<=Vw;
XbG_H178<=Vw;
XbG_H179<=Vw;
XbG_H18<=Vw;
XbG_H180<=Vw;
XbG_H181<=Vw;
XbG_H182<=Vw;
XbG_H183<=Vw;
XbG_H184<=Vw;
XbG_H185<=Vw;
XbG_H186<=Vw;
XbG_H187<=Vw;
XbG_H188<=Vw;
XbG_H189<=Vw;
XbG_H19<=Vw;
XbG_H190<=Vw;
XbG_H191<=Vw;
XbG_H192<=Vw;
XbG_H193<=Vw;
XbG_H194<=Vw;
XbG_H195<=Vw;
XbG_H196<=Vw;
XbG_H197<=Vw;
XbG_H198<=Vw;
XbG_H199<=Vw;
XbG_H2<=Vw;
XbG_H20<=Vw;
XbG_H200<=Vw;
XbG_H201<=Vw;
XbG_H202<=Vw;
XbG_H203<=Vw;
XbG_H204<=Vw;
XbG_H205<=Vw;
XbG_H206<=Vw;
XbG_H207<=Vw;
XbG_H208<=Vw;
XbG_H209<=Vw;
XbG_H21<=Vw;
XbG_H210<=Vw;
XbG_H211<=Vw;
XbG_H212<=Vw;
XbG_H213<=Vw;
XbG_H214<=Vw;
XbG_H215<=Vw;
XbG_H216<=Vw;
XbG_H217<=Vw;
XbG_H218<=Vw;
XbG_H219<=Vw;
XbG_H22<=Vw;
XbG_H220<=Vw;
XbG_H221<=Vw;
XbG_H222<=Vw;
XbG_H223<=Vw;
XbG_H224<=Vw;
XbG_H225<=Vw;
XbG_H226<=Vw;
XbG_H227<=Vw;
XbG_H228<=Vw;
XbG_H229<=Vw;
XbG_H23<=Vw;
XbG_H230<=Vw;
XbG_H231<=Vw;
XbG_H232<=Vw;
XbG_H233<=Vw;
XbG_H234<=Vw;
XbG_H235<=Vw;
XbG_H236<=Vw;
XbG_H237<=Vw;
XbG_H238<=Vw;
XbG_H239<=Vw;
XbG_H24<=Vw;
XbG_H240<=Vw;
XbG_H241<=Vw;
XbG_H242<=Vw;
XbG_H243<=Vw;
XbG_H244<=Vw;
XbG_H245<=Vw;
XbG_H246<=Vw;
XbG_H247<=Vw;
XbG_H248<=Vw;
XbG_H249<=Vw;
XbG_H25<=Vw;
XbG_H250<=Vw;
XbG_H251<=Vw;
XbG_H252<=Vw;
XbG_H253<=Vw;
XbG_H254<=Vw;
XbG_H255<=Vw;
XbG_H256<=Vw;
XbG_H257<=Vw;
XbG_H258<=Vw;
XbG_H259<=Vw;
XbG_H26<=Vw;
XbG_H260<=Vw;
XbG_H261<=Vw;
XbG_H262<=Vw;
XbG_H263<=Vw;
XbG_H264<=Vw;
XbG_H265<=Vw;
XbG_H266<=Vw;
XbG_H267<=Vw;
XbG_H268<=Vw;
XbG_H269<=Vw;
XbG_H27<=Vw;
XbG_H270<=Vw;
XbG_H271<=Vw;
XbG_H272<=Vw;
XbG_H273<=Vw;
XbG_H274<=Vw;
XbG_H275<=Vw;
XbG_H276<=Vw;
XbG_H277<=Vw;
XbG_H278<=Vw;
XbG_H279<=Vw;
XbG_H28<=Vw;
XbG_H280<=Vw;
XbG_H281<=Vw;
XbG_H282<=Vw;
XbG_H283<=Vw;
XbG_H284<=Vw;
XbG_H285<=Vw;
XbG_H286<=Vw;
XbG_H287<=Vw;
XbG_H288<=Vw;
XbG_H289<=Vw;
XbG_H29<=Vw;
XbG_H290<=Vw;
XbG_H291<=Vw;
XbG_H292<=Vw;
XbG_H293<=Vw;
XbG_H294<=Vw;
XbG_H295<=Vw;
XbG_H296<=Vw;
XbG_H297<=Vw;
XbG_H298<=Vw;
XbG_H299<=Vw;
XbG_H3<=Vw;
XbG_H30<=Vw;
XbG_H300<=Vw;
XbG_H301<=Vw;
XbG_H302<=Vw;
XbG_H303<=Vw;
XbG_H304<=Vw;
XbG_H305<=Vw;
XbG_H306<=Vw;
XbG_H307<=Vw;
XbG_H308<=Vw;
XbG_H309<=Vw;
XbG_H31<=Vw;
XbG_H310<=Vw;
XbG_H311<=Vw;
XbG_H312<=Vw;
XbG_H313<=Vw;
XbG_H314<=Vw;
XbG_H315<=Vw;
XbG_H316<=Vw;
XbG_H317<=Vw;
XbG_H318<=Vw;
XbG_H319<=Vw;
XbG_H32<=Vw;
XbG_H320<=Vw;
XbG_H321<=Vw;
XbG_H322<=Vw;
XbG_H323<=Vw;
XbG_H324<=Vw;
XbG_H325<=Vw;
XbG_H326<=Vw;
XbG_H327<=Vw;
XbG_H328<=Vw;
XbG_H329<=Vw;
XbG_H33<=Vw;
XbG_H330<=Vw;
XbG_H331<=Vw;
XbG_H332<=Vw;
XbG_H333<=Vw;
XbG_H334<=Vw;
XbG_H335<=Vw;
XbG_H336<=Vw;
XbG_H337<=Vw;
XbG_H338<=Vw;
XbG_H339<=Vw;
XbG_H34<=Vw;
XbG_H340<=Vw;
XbG_H341<=Vw;
XbG_H342<=Vw;
XbG_H343<=Vw;
XbG_H344<=Vw;
XbG_H345<=Vw;
XbG_H346<=Vw;
XbG_H347<=Vw;
XbG_H348<=Vw;
XbG_H349<=Vw;
XbG_H35<=Vw;
XbG_H350<=Vw;
XbG_H351<=Vw;
XbG_H352<=Vw;
XbG_H353<=Vw;
XbG_H354<=Vw;
XbG_H355<=Vw;
XbG_H356<=Vw;
XbG_H357<=Vw;
XbG_H358<=Vw;
XbG_H359<=Vw;
XbG_H36<=Vw;
XbG_H360<=Vw;
XbG_H361<=Vw;
XbG_H362<=Vw;
XbG_H363<=Vw;
XbG_H364<=Vw;
XbG_H365<=Vw;
XbG_H366<=Vw;
XbG_H367<=Vw;
XbG_H368<=Vw;
XbG_H369<=Vw;
XbG_H37<=Vw;
XbG_H370<=Vw;
XbG_H371<=Vw;
XbG_H372<=Vw;
XbG_H373<=Vw;
XbG_H374<=Vw;
XbG_H375<=Vw;
XbG_H376<=Vw;
XbG_H377<=Vw;
XbG_H378<=Vw;
XbG_H379<=Vw;
XbG_H38<=Vw;
XbG_H380<=Vw;
XbG_H381<=Vw;
XbG_H382<=Vw;
XbG_H383<=Vw;
XbG_H384<=Vw;
XbG_H385<=Vw;
XbG_H386<=Vw;
XbG_H387<=Vw;
XbG_H388<=Vw;
XbG_H389<=Vw;
XbG_H39<=Vw;
XbG_H390<=Vw;
XbG_H391<=Vw;
XbG_H392<=Vw;
XbG_H393<=Vw;
XbG_H394<=Vw;
XbG_H395<=Vw;
XbG_H396<=Vw;
XbG_H397<=Vw;
XbG_H398<=Vw;
XbG_H399<=Vw;
XbG_H4<=Vw;
XbG_H40<=Vw;
XbG_H400<=Vw;
XbG_H401<=Vw;
XbG_H402<=Vw;
XbG_H403<=Vw;
XbG_H404<=Vw;
XbG_H405<=Vw;
XbG_H406<=Vw;
XbG_H407<=Vw;
XbG_H408<=Vw;
XbG_H409<=Vw;
XbG_H41<=Vw;
XbG_H410<=Vw;
XbG_H411<=Vw;
XbG_H412<=Vw;
XbG_H413<=Vw;
XbG_H414<=Vw;
XbG_H415<=Vw;
XbG_H416<=Vw;
XbG_H417<=Vw;
XbG_H418<=Vw;
XbG_H419<=Vw;
XbG_H42<=Vw;
XbG_H420<=Vw;
XbG_H421<=Vw;
XbG_H422<=Vw;
XbG_H423<=Vw;
XbG_H424<=Vw;
XbG_H425<=Vw;
XbG_H426<=Vw;
XbG_H427<=Vw;
XbG_H428<=Vw;
XbG_H429<=Vw;
XbG_H43<=Vw;
XbG_H430<=Vw;
XbG_H431<=Vw;
XbG_H432<=Vw;
XbG_H433<=Vw;
XbG_H434<=Vw;
XbG_H435<=Vw;
XbG_H436<=Vw;
XbG_H437<=Vw;
XbG_H438<=Vw;
XbG_H439<=Vw;
XbG_H44<=Vw;
XbG_H440<=Vw;
XbG_H441<=Vw;
XbG_H442<=Vw;
XbG_H443<=Vw;
XbG_H444<=Vw;
XbG_H445<=Vw;
XbG_H446<=Vw;
XbG_H447<=Vw;
XbG_H448<=Vw;
XbG_H449<=Vw;
XbG_H45<=Vw;
XbG_H450<=Vw;
XbG_H451<=Vw;
XbG_H452<=Vw;
XbG_H453<=Vw;
XbG_H454<=Vw;
XbG_H455<=Vw;
XbG_H456<=Vw;
XbG_H457<=Vw;
XbG_H458<=Vw;
XbG_H459<=Vw;
XbG_H46<=Vw;
XbG_H460<=Vw;
XbG_H461<=Vw;
XbG_H462<=Vw;
XbG_H463<=Vw;
XbG_H464<=Vw;
XbG_H465<=Vw;
XbG_H466<=Vw;
XbG_H467<=Vw;
XbG_H468<=Vw;
XbG_H469<=Vw;
XbG_H47<=Vw;
XbG_H470<=Vw;
XbG_H471<=Vw;
XbG_H472<=Vw;
XbG_H473<=Vw;
XbG_H474<=Vw;
XbG_H475<=Vw;
XbG_H476<=Vw;
XbG_H477<=Vw;
XbG_H478<=Vw;
XbG_H479<=Vw;
XbG_H48<=Vw;
XbG_H480<=Vw;
XbG_H481<=Vw;
XbG_H482<=Vw;
XbG_H483<=Vw;
XbG_H484<=Vw;
XbG_H485<=Vw;
XbG_H486<=Vw;
XbG_H487<=Vw;
XbG_H488<=Vw;
XbG_H489<=Vw;
XbG_H49<=Vw;
XbG_H490<=Vw;
XbG_H491<=Vw;
XbG_H492<=Vw;
XbG_H493<=Vw;
XbG_H494<=Vw;
XbG_H495<=Vw;
XbG_H496<=Vw;
XbG_H497<=Vw;
XbG_H498<=Vw;
XbG_H499<=Vw;
XbG_H5<=Vw;
XbG_H50<=Vw;
XbG_H500<=Vw;
XbG_H501<=Vw;
XbG_H502<=Vw;
XbG_H503<=Vw;
XbG_H504<=Vw;
XbG_H505<=Vw;
XbG_H506<=Vw;
XbG_H507<=Vw;
XbG_H508<=Vw;
XbG_H509<=Vw;
XbG_H51<=Vw;
XbG_H510<=Vw;
XbG_H511<=Vw;
XbG_H512<=Vw;
XbG_H513<=Vw;
XbG_H514<=Vw;
XbG_H515<=Vw;
XbG_H516<=Vw;
XbG_H517<=Vw;
XbG_H518<=Vw;
XbG_H519<=Vw;
XbG_H52<=Vw;
XbG_H520<=Vw;
XbG_H521<=Vw;
XbG_H522<=Vw;
XbG_H523<=Vw;
XbG_H524<=Vw;
XbG_H525<=Vw;
XbG_H526<=Vw;
XbG_H527<=Vw;
XbG_H528<=Vw;
XbG_H529<=Vw;
XbG_H53<=Vw;
XbG_H530<=Vw;
XbG_H531<=Vw;
XbG_H532<=Vw;
XbG_H533<=Vw;
XbG_H534<=Vw;
XbG_H535<=Vw;
XbG_H536<=Vw;
XbG_H537<=Vw;
XbG_H538<=Vw;
XbG_H539<=Vw;
XbG_H54<=Vw;
XbG_H540<=Vw;
XbG_H541<=Vw;
XbG_H542<=Vw;
XbG_H543<=Vw;
XbG_H544<=Vw;
XbG_H545<=Vw;
XbG_H546<=Vw;
XbG_H547<=Vw;
XbG_H548<=Vw;
XbG_H549<=Vw;
XbG_H55<=Vw;
XbG_H550<=Vw;
XbG_H551<=Vw;
XbG_H552<=Vw;
XbG_H553<=Vw;
XbG_H554<=Vw;
XbG_H555<=Vw;
XbG_H556<=Vw;
XbG_H557<=Vw;
XbG_H558<=Vw;
XbG_H559<=Vw;
XbG_H56<=Vw;
XbG_H560<=Vw;
XbG_H561<=Vw;
XbG_H562<=Vw;
XbG_H563<=Vw;
XbG_H564<=Vw;
XbG_H565<=Vw;
XbG_H566<=Vw;
XbG_H567<=Vw;
XbG_H568<=Vw;
XbG_H569<=Vw;
XbG_H57<=Vw;
XbG_H570<=Vw;
XbG_H571<=Vw;
XbG_H572<=Vw;
XbG_H573<=Vw;
XbG_H574<=Vw;
XbG_H575<=Vw;
XbG_H576<=Vw;
XbG_H577<=Vw;
XbG_H578<=Vw;
XbG_H579<=Vw;
XbG_H58<=Vw;
XbG_H580<=Vw;
XbG_H581<=Vw;
XbG_H582<=Vw;
XbG_H583<=Vw;
XbG_H584<=Vw;
XbG_H585<=Vw;
XbG_H586<=Vw;
XbG_H587<=Vw;
XbG_H588<=Vw;
XbG_H589<=Vw;
XbG_H59<=Vw;
XbG_H590<=Vw;
XbG_H591<=Vw;
XbG_H592<=Vw;
XbG_H593<=Vw;
XbG_H594<=Vw;
XbG_H595<=Vw;
XbG_H596<=Vw;
XbG_H597<=Vw;
XbG_H598<=Vw;
XbG_H599<=Vw;
XbG_H6<=Vw;
XbG_H60<=Vw;
XbG_H600<=Vw;
XbG_H601<=Vw;
XbG_H602<=Vw;
XbG_H603<=Vw;
XbG_H604<=Vw;
XbG_H605<=Vw;
XbG_H606<=Vw;
XbG_H607<=Vw;
XbG_H608<=Vw;
XbG_H609<=Vw;
XbG_H61<=Vw;
XbG_H610<=Vw;
XbG_H611<=Vw;
XbG_H612<=Vw;
XbG_H613<=Vw;
XbG_H614<=Vw;
XbG_H615<=Vw;
XbG_H616<=Vw;
XbG_H617<=Vw;
XbG_H618<=Vw;
XbG_H619<=Vw;
XbG_H62<=Vw;
XbG_H620<=Vw;
XbG_H621<=Vw;
XbG_H622<=Vw;
XbG_H623<=Vw;
XbG_H624<=Vw;
XbG_H625<=Vw;
XbG_H626<=Vw;
XbG_H627<=Vw;
XbG_H628<=Vw;
XbG_H629<=Vw;
XbG_H63<=Vw;
XbG_H630<=Vw;
XbG_H631<=Vw;
XbG_H632<=Vw;
XbG_H633<=Vw;
XbG_H634<=Vw;
XbG_H635<=Vw;
XbG_H636<=Vw;
XbG_H637<=Vw;
XbG_H638<=Vw;
XbG_H639<=Vw;
XbG_H64<=Vw;
XbG_H640<=Vw;
XbG_H641<=Vw;
XbG_H642<=Vw;
XbG_H643<=Vw;
XbG_H644<=Vw;
XbG_H645<=Vw;
XbG_H646<=Vw;
XbG_H647<=Vw;
XbG_H648<=Vw;
XbG_H649<=Vw;
XbG_H65<=Vw;
XbG_H650<=Vw;
XbG_H651<=Vw;
XbG_H652<=Vw;
XbG_H653<=Vw;
XbG_H654<=Vw;
XbG_H655<=Vw;
XbG_H656<=Vw;
XbG_H657<=Vw;
XbG_H658<=Vw;
XbG_H659<=Vw;
XbG_H66<=Vw;
XbG_H660<=Vw;
XbG_H661<=Vw;
XbG_H662<=Vw;
XbG_H663<=Vw;
XbG_H664<=Vw;
XbG_H665<=Vw;
XbG_H666<=Vw;
XbG_H667<=Vw;
XbG_H668<=Vw;
XbG_H669<=Vw;
XbG_H67<=Vw;
XbG_H670<=Vw;
XbG_H671<=Vw;
XbG_H672<=Vw;
XbG_H673<=Vw;
XbG_H674<=Vw;
XbG_H675<=Vw;
XbG_H676<=Vw;
XbG_H677<=Vw;
XbG_H678<=Vw;
XbG_H679<=Vw;
XbG_H68<=Vw;
XbG_H680<=Vw;
XbG_H681<=Vw;
XbG_H682<=Vw;
XbG_H683<=Vw;
XbG_H684<=Vw;
XbG_H685<=Vw;
XbG_H686<=Vw;
XbG_H687<=Vw;
XbG_H688<=Vw;
XbG_H689<=Vw;
XbG_H69<=Vw;
XbG_H690<=Vw;
XbG_H691<=Vw;
XbG_H692<=Vw;
XbG_H693<=Vw;
XbG_H694<=Vw;
XbG_H695<=Vw;
XbG_H696<=Vw;
XbG_H697<=Vw;
XbG_H698<=Vw;
XbG_H699<=Vw;
XbG_H7<=Vw;
XbG_H70<=Vw;
XbG_H700<=Vw;
XbG_H701<=Vw;
XbG_H702<=Vw;
XbG_H703<=Vw;
XbG_H704<=Vw;
XbG_H705<=Vw;
XbG_H706<=Vw;
XbG_H707<=Vw;
XbG_H708<=Vw;
XbG_H709<=Vw;
XbG_H71<=Vw;
XbG_H710<=Vw;
XbG_H711<=Vw;
XbG_H712<=Vw;
XbG_H713<=Vw;
XbG_H714<=Vw;
XbG_H715<=Vw;
XbG_H716<=Vw;
XbG_H717<=Vw;
XbG_H718<=Vw;
XbG_H719<=Vw;
XbG_H72<=Vw;
XbG_H720<=Vw;
XbG_H721<=Vw;
XbG_H722<=Vw;
XbG_H723<=Vw;
XbG_H724<=Vw;
XbG_H725<=Vw;
XbG_H726<=Vw;
XbG_H727<=Vw;
XbG_H728<=Vw;
XbG_H729<=Vw;
XbG_H73<=Vw;
XbG_H730<=Vw;
XbG_H731<=Vw;
XbG_H732<=Vw;
XbG_H733<=Vw;
XbG_H734<=Vw;
XbG_H735<=Vw;
XbG_H74<=Vw;
XbG_H75<=Vw;
XbG_H76<=Vw;
XbG_H77<=Vw;
XbG_H78<=Vw;
XbG_H79<=Vw;
XbG_H8<=Vw;
XbG_H80<=Vw;
XbG_H81<=Vw;
XbG_H82<=Vw;
XbG_H83<=Vw;
XbG_H84<=Vw;
XbG_H85<=Vw;
XbG_H86<=Vw;
XbG_H87<=Vw;
XbG_H88<=Vw;
XbG_H89<=Vw;
XbG_H9<=Vw;
XbG_H90<=Vw;
XbG_H91<=Vw;
XbG_H92<=Vw;
XbG_H93<=Vw;
XbG_H94<=Vw;
XbG_H95<=Vw;
XbG_H96<=Vw;
XbG_H97<=Vw;
XbG_H98<=Vw;
XbG_H99<=Vw;
XbG_V0<=zero;
XbG_V1<=zero;
XbG_V10<=zero;
XbG_V100<=zero;
XbG_V101<=zero;
XbG_V102<=zero;
XbG_V103<=zero;
XbG_V104<=zero;
XbG_V105<=zero;
XbG_V106<=zero;
XbG_V107<=zero;
XbG_V108<=zero;
XbG_V109<=zero;
XbG_V11<=zero;
XbG_V110<=zero;
XbG_V111<=zero;
XbG_V112<=zero;
XbG_V113<=zero;
XbG_V114<=zero;
XbG_V115<=zero;
XbG_V116<=zero;
XbG_V117<=zero;
XbG_V118<=zero;
XbG_V119<=zero;
XbG_V12<=zero;
XbG_V120<=zero;
XbG_V121<=zero;
XbG_V122<=zero;
XbG_V123<=zero;
XbG_V124<=zero;
XbG_V125<=zero;
XbG_V126<=zero;
XbG_V127<=zero;
XbG_V128<=zero;
XbG_V129<=zero;
XbG_V13<=zero;
XbG_V130<=zero;
XbG_V131<=zero;
XbG_V132<=zero;
XbG_V133<=zero;
XbG_V134<=zero;
XbG_V135<=zero;
XbG_V136<=zero;
XbG_V137<=zero;
XbG_V138<=zero;
XbG_V139<=zero;
XbG_V14<=zero;
XbG_V140<=zero;
XbG_V141<=zero;
XbG_V142<=zero;
XbG_V143<=zero;
XbG_V144<=zero;
XbG_V145<=zero;
XbG_V146<=zero;
XbG_V147<=zero;
XbG_V148<=zero;
XbG_V149<=zero;
XbG_V15<=zero;
XbG_V150<=zero;
XbG_V151<=zero;
XbG_V152<=zero;
XbG_V153<=zero;
XbG_V154<=zero;
XbG_V155<=zero;
XbG_V156<=zero;
XbG_V157<=zero;
XbG_V158<=zero;
XbG_V159<=zero;
XbG_V16<=zero;
XbG_V160<=zero;
XbG_V161<=zero;
XbG_V162<=zero;
XbG_V163<=zero;
XbG_V164<=zero;
XbG_V165<=zero;
XbG_V166<=zero;
XbG_V167<=zero;
XbG_V168<=zero;
XbG_V169<=zero;
XbG_V17<=zero;
XbG_V170<=zero;
XbG_V171<=zero;
XbG_V172<=zero;
XbG_V173<=zero;
XbG_V174<=zero;
XbG_V175<=zero;
XbG_V176<=zero;
XbG_V177<=zero;
XbG_V178<=zero;
XbG_V179<=zero;
XbG_V18<=zero;
XbG_V180<=zero;
XbG_V181<=zero;
XbG_V182<=zero;
XbG_V183<=zero;
XbG_V184<=zero;
XbG_V185<=zero;
XbG_V186<=zero;
XbG_V187<=zero;
XbG_V188<=zero;
XbG_V189<=zero;
XbG_V19<=zero;
XbG_V2<=zero;
XbG_V20<=zero;
XbG_V21<=zero;
XbG_V22<=zero;
XbG_V23<=zero;
XbG_V24<=zero;
XbG_V25<=zero;
XbG_V26<=zero;
XbG_V27<=zero;
XbG_V28<=zero;
XbG_V29<=zero;
XbG_V3<=zero;
XbG_V30<=zero;
XbG_V31<=zero;
XbG_V32<=zero;
XbG_V33<=zero;
XbG_V34<=zero;
XbG_V35<=zero;
XbG_V36<=zero;
XbG_V37<=zero;
XbG_V38<=zero;
XbG_V39<=zero;
XbG_V4<=zero;
XbG_V40<=zero;
XbG_V41<=zero;
XbG_V42<=zero;
XbG_V43<=zero;
XbG_V44<=zero;
XbG_V45<=zero;
XbG_V46<=zero;
XbG_V47<=zero;
XbG_V48<=zero;
XbG_V49<=zero;
XbG_V5<=zero;
XbG_V50<=zero;
XbG_V51<=zero;
XbG_V52<=zero;
XbG_V53<=zero;
XbG_V54<=zero;
XbG_V55<=zero;
XbG_V56<=zero;
XbG_V57<=zero;
XbG_V58<=zero;
XbG_V59<=zero;
XbG_V6<=zero;
XbG_V60<=zero;
XbG_V61<=zero;
XbG_V62<=zero;
XbG_V63<=zero;
XbG_V64<=zero;
XbG_V65<=zero;
XbG_V66<=zero;
XbG_V67<=zero;
XbG_V68<=zero;
XbG_V69<=zero;
XbG_V7<=zero;
XbG_V70<=zero;
XbG_V71<=zero;
XbG_V72<=zero;
XbG_V73<=zero;
XbG_V74<=zero;
XbG_V75<=zero;
XbG_V76<=zero;
XbG_V77<=zero;
XbG_V78<=zero;
XbG_V79<=zero;
XbG_V8<=zero;
XbG_V80<=zero;
XbG_V81<=zero;
XbG_V82<=zero;
XbG_V83<=zero;
XbG_V84<=zero;
XbG_V85<=zero;
XbG_V86<=zero;
XbG_V87<=zero;
XbG_V88<=zero;
XbG_V89<=zero;
XbG_V9<=zero;
XbG_V90<=zero;
XbG_V91<=zero;
XbG_V92<=zero;
XbG_V93<=zero;
XbG_V94<=zero;
XbG_V95<=zero;
XbG_V96<=zero;
XbG_V97<=zero;
XbG_V98<=zero;
XbG_V99<=zero;

else

XbG_H0<=Vw;
XbG_H1<=Vw;
XbG_H10<=Vw;
XbG_H100<=Vw;
XbG_H101<=Vw;
XbG_H102<=Vw;
XbG_H103<=Vw;
XbG_H104<=Vw;
XbG_H105<=Vw;
XbG_H106<=Vw;
XbG_H107<=Vw;
XbG_H108<=Vw;
XbG_H109<=Vw;
XbG_H11<=Vw;
XbG_H110<=Vw;
XbG_H111<=Vw;
XbG_H112<=Vw;
XbG_H113<=Vw;
XbG_H114<=Vw;
XbG_H115<=Vw;
XbG_H116<=Vw;
XbG_H117<=Vw;
XbG_H118<=Vw;
XbG_H119<=Vw;
XbG_H12<=Vw;
XbG_H120<=Vw;
XbG_H121<=Vw;
XbG_H122<=Vw;
XbG_H123<=Vw;
XbG_H124<=Vw;
XbG_H125<=Vw;
XbG_H126<=Vw;
XbG_H127<=Vw;
XbG_H128<=Vw;
XbG_H129<=Vw;
XbG_H13<=Vw;
XbG_H130<=Vw;
XbG_H131<=Vw;
XbG_H132<=Vw;
XbG_H133<=Vw;
XbG_H134<=Vw;
XbG_H135<=Vw;
XbG_H136<=Vw;
XbG_H137<=Vw;
XbG_H138<=Vw;
XbG_H139<=Vw;
XbG_H14<=Vw;
XbG_H140<=Vw;
XbG_H141<=Vw;
XbG_H142<=Vw;
XbG_H143<=Vw;
XbG_H144<=Vw;
XbG_H145<=Vw;
XbG_H146<=Vw;
XbG_H147<=Vw;
XbG_H148<=Vw;
XbG_H149<=Vw;
XbG_H15<=Vw;
XbG_H150<=Vw;
XbG_H151<=Vw;
XbG_H152<=Vw;
XbG_H153<=Vw;
XbG_H154<=Vw;
XbG_H155<=Vw;
XbG_H156<=Vw;
XbG_H157<=Vw;
XbG_H158<=Vw;
XbG_H159<=Vw;
XbG_H16<=Vw;
XbG_H160<=Vw;
XbG_H161<=Vw;
XbG_H162<=Vw;
XbG_H163<=Vw;
XbG_H164<=Vw;
XbG_H165<=Vw;
XbG_H166<=Vw;
XbG_H167<=Vw;
XbG_H168<=Vw;
XbG_H169<=Vw;
XbG_H17<=Vw;
XbG_H170<=Vw;
XbG_H171<=Vw;
XbG_H172<=Vw;
XbG_H173<=Vw;
XbG_H174<=Vw;
XbG_H175<=Vw;
XbG_H176<=Vw;
XbG_H177<=Vw;
XbG_H178<=Vw;
XbG_H179<=Vw;
XbG_H18<=Vw;
XbG_H180<=Vw;
XbG_H181<=Vw;
XbG_H182<=Vw;
XbG_H183<=Vw;
XbG_H184<=Vw;
XbG_H185<=Vw;
XbG_H186<=Vw;
XbG_H187<=Vw;
XbG_H188<=Vw;
XbG_H189<=Vw;
XbG_H19<=Vw;
XbG_H190<=Vw;
XbG_H191<=Vw;
XbG_H192<=Vw;
XbG_H193<=Vw;
XbG_H194<=Vw;
XbG_H195<=Vw;
XbG_H196<=Vw;
XbG_H197<=Vw;
XbG_H198<=Vw;
XbG_H199<=Vw;
XbG_H2<=Vw;
XbG_H20<=Vw;
XbG_H200<=Vw;
XbG_H201<=Vw;
XbG_H202<=Vw;
XbG_H203<=Vw;
XbG_H204<=Vw;
XbG_H205<=Vw;
XbG_H206<=Vw;
XbG_H207<=Vw;
XbG_H208<=Vw;
XbG_H209<=Vw;
XbG_H21<=Vw;
XbG_H210<=Vw;
XbG_H211<=Vw;
XbG_H212<=Vw;
XbG_H213<=Vw;
XbG_H214<=Vw;
XbG_H215<=Vw;
XbG_H216<=Vw;
XbG_H217<=Vw;
XbG_H218<=Vw;
XbG_H219<=Vw;
XbG_H22<=Vw;
XbG_H220<=Vw;
XbG_H221<=Vw;
XbG_H222<=Vw;
XbG_H223<=Vw;
XbG_H224<=Vw;
XbG_H225<=Vw;
XbG_H226<=Vw;
XbG_H227<=Vw;
XbG_H228<=Vw;
XbG_H229<=Vw;
XbG_H23<=Vw;
XbG_H230<=Vw;
XbG_H231<=Vw;
XbG_H232<=Vw;
XbG_H233<=Vw;
XbG_H234<=Vw;
XbG_H235<=Vw;
XbG_H236<=Vw;
XbG_H237<=Vw;
XbG_H238<=Vw;
XbG_H239<=Vw;
XbG_H24<=Vw;
XbG_H240<=Vw;
XbG_H241<=Vw;
XbG_H242<=Vw;
XbG_H243<=Vw;
XbG_H244<=Vw;
XbG_H245<=Vw;
XbG_H246<=Vw;
XbG_H247<=Vw;
XbG_H248<=Vw;
XbG_H249<=Vw;
XbG_H25<=Vw;
XbG_H250<=Vw;
XbG_H251<=Vw;
XbG_H252<=Vw;
XbG_H253<=Vw;
XbG_H254<=Vw;
XbG_H255<=Vw;
XbG_H256<=Vw;
XbG_H257<=Vw;
XbG_H258<=Vw;
XbG_H259<=Vw;
XbG_H26<=Vw;
XbG_H260<=Vw;
XbG_H261<=Vw;
XbG_H262<=Vw;
XbG_H263<=Vw;
XbG_H264<=Vw;
XbG_H265<=Vw;
XbG_H266<=Vw;
XbG_H267<=Vw;
XbG_H268<=Vw;
XbG_H269<=Vw;
XbG_H27<=Vw;
XbG_H270<=Vw;
XbG_H271<=Vw;
XbG_H272<=Vw;
XbG_H273<=Vw;
XbG_H274<=Vw;
XbG_H275<=Vw;
XbG_H276<=Vw;
XbG_H277<=Vw;
XbG_H278<=Vw;
XbG_H279<=Vw;
XbG_H28<=Vw;
XbG_H280<=Vw;
XbG_H281<=Vw;
XbG_H282<=Vw;
XbG_H283<=Vw;
XbG_H284<=Vw;
XbG_H285<=Vw;
XbG_H286<=Vw;
XbG_H287<=Vw;
XbG_H288<=Vw;
XbG_H289<=Vw;
XbG_H29<=Vw;
XbG_H290<=Vw;
XbG_H291<=Vw;
XbG_H292<=Vw;
XbG_H293<=Vw;
XbG_H294<=Vw;
XbG_H295<=Vw;
XbG_H296<=Vw;
XbG_H297<=Vw;
XbG_H298<=Vw;
XbG_H299<=Vw;
XbG_H3<=Vw;
XbG_H30<=Vw;
XbG_H300<=Vw;
XbG_H301<=Vw;
XbG_H302<=Vw;
XbG_H303<=Vw;
XbG_H304<=Vw;
XbG_H305<=Vw;
XbG_H306<=Vw;
XbG_H307<=Vw;
XbG_H308<=Vw;
XbG_H309<=Vw;
XbG_H31<=Vw;
XbG_H310<=Vw;
XbG_H311<=Vw;
XbG_H312<=Vw;
XbG_H313<=Vw;
XbG_H314<=Vw;
XbG_H315<=Vw;
XbG_H316<=Vw;
XbG_H317<=Vw;
XbG_H318<=Vw;
XbG_H319<=Vw;
XbG_H32<=Vw;
XbG_H320<=Vw;
XbG_H321<=Vw;
XbG_H322<=Vw;
XbG_H323<=Vw;
XbG_H324<=Vw;
XbG_H325<=Vw;
XbG_H326<=Vw;
XbG_H327<=Vw;
XbG_H328<=Vw;
XbG_H329<=Vw;
XbG_H33<=Vw;
XbG_H330<=Vw;
XbG_H331<=Vw;
XbG_H332<=Vw;
XbG_H333<=Vw;
XbG_H334<=Vw;
XbG_H335<=Vw;
XbG_H336<=Vw;
XbG_H337<=Vw;
XbG_H338<=Vw;
XbG_H339<=Vw;
XbG_H34<=Vw;
XbG_H340<=Vw;
XbG_H341<=Vw;
XbG_H342<=Vw;
XbG_H343<=Vw;
XbG_H344<=Vw;
XbG_H345<=Vw;
XbG_H346<=Vw;
XbG_H347<=Vw;
XbG_H348<=Vw;
XbG_H349<=Vw;
XbG_H35<=Vw;
XbG_H350<=Vw;
XbG_H351<=Vw;
XbG_H352<=Vw;
XbG_H353<=Vw;
XbG_H354<=Vw;
XbG_H355<=Vw;
XbG_H356<=Vw;
XbG_H357<=Vw;
XbG_H358<=Vw;
XbG_H359<=Vw;
XbG_H36<=Vw;
XbG_H360<=Vw;
XbG_H361<=Vw;
XbG_H362<=Vw;
XbG_H363<=Vw;
XbG_H364<=Vw;
XbG_H365<=Vw;
XbG_H366<=Vw;
XbG_H367<=Vw;
XbG_H368<=Vw;
XbG_H369<=Vw;
XbG_H37<=Vw;
XbG_H370<=Vw;
XbG_H371<=Vw;
XbG_H372<=Vw;
XbG_H373<=Vw;
XbG_H374<=Vw;
XbG_H375<=Vw;
XbG_H376<=Vw;
XbG_H377<=Vw;
XbG_H378<=Vw;
XbG_H379<=Vw;
XbG_H38<=Vw;
XbG_H380<=Vw;
XbG_H381<=Vw;
XbG_H382<=Vw;
XbG_H383<=Vw;
XbG_H384<=Vw;
XbG_H385<=Vw;
XbG_H386<=Vw;
XbG_H387<=Vw;
XbG_H388<=Vw;
XbG_H389<=Vw;
XbG_H39<=Vw;
XbG_H390<=Vw;
XbG_H391<=Vw;
XbG_H392<=Vw;
XbG_H393<=Vw;
XbG_H394<=Vw;
XbG_H395<=Vw;
XbG_H396<=Vw;
XbG_H397<=Vw;
XbG_H398<=Vw;
XbG_H399<=Vw;
XbG_H4<=Vw;
XbG_H40<=Vw;
XbG_H400<=Vw;
XbG_H401<=Vw;
XbG_H402<=Vw;
XbG_H403<=Vw;
XbG_H404<=Vw;
XbG_H405<=Vw;
XbG_H406<=Vw;
XbG_H407<=Vw;
XbG_H408<=Vw;
XbG_H409<=Vw;
XbG_H41<=Vw;
XbG_H410<=Vw;
XbG_H411<=Vw;
XbG_H412<=Vw;
XbG_H413<=Vw;
XbG_H414<=Vw;
XbG_H415<=Vw;
XbG_H416<=Vw;
XbG_H417<=Vw;
XbG_H418<=Vw;
XbG_H419<=Vw;
XbG_H42<=Vw;
XbG_H420<=Vw;
XbG_H421<=Vw;
XbG_H422<=Vw;
XbG_H423<=Vw;
XbG_H424<=Vw;
XbG_H425<=Vw;
XbG_H426<=Vw;
XbG_H427<=Vw;
XbG_H428<=Vw;
XbG_H429<=Vw;
XbG_H43<=Vw;
XbG_H430<=Vw;
XbG_H431<=Vw;
XbG_H432<=Vw;
XbG_H433<=Vw;
XbG_H434<=Vw;
XbG_H435<=Vw;
XbG_H436<=Vw;
XbG_H437<=Vw;
XbG_H438<=Vw;
XbG_H439<=Vw;
XbG_H44<=Vw;
XbG_H440<=Vw;
XbG_H441<=Vw;
XbG_H442<=Vw;
XbG_H443<=Vw;
XbG_H444<=Vw;
XbG_H445<=Vw;
XbG_H446<=Vw;
XbG_H447<=Vw;
XbG_H448<=Vw;
XbG_H449<=Vw;
XbG_H45<=Vw;
XbG_H450<=Vw;
XbG_H451<=Vw;
XbG_H452<=Vw;
XbG_H453<=Vw;
XbG_H454<=Vw;
XbG_H455<=Vw;
XbG_H456<=Vw;
XbG_H457<=Vw;
XbG_H458<=Vw;
XbG_H459<=Vw;
XbG_H46<=Vw;
XbG_H460<=Vw;
XbG_H461<=Vw;
XbG_H462<=Vw;
XbG_H463<=Vw;
XbG_H464<=Vw;
XbG_H465<=Vw;
XbG_H466<=Vw;
XbG_H467<=Vw;
XbG_H468<=Vw;
XbG_H469<=Vw;
XbG_H47<=Vw;
XbG_H470<=Vw;
XbG_H471<=Vw;
XbG_H472<=Vw;
XbG_H473<=Vw;
XbG_H474<=Vw;
XbG_H475<=Vw;
XbG_H476<=Vw;
XbG_H477<=Vw;
XbG_H478<=Vw;
XbG_H479<=Vw;
XbG_H48<=Vw;
XbG_H480<=Vw;
XbG_H481<=Vw;
XbG_H482<=Vw;
XbG_H483<=Vw;
XbG_H484<=Vw;
XbG_H485<=Vw;
XbG_H486<=Vw;
XbG_H487<=Vw;
XbG_H488<=Vw;
XbG_H489<=Vw;
XbG_H49<=Vw;
XbG_H490<=Vw;
XbG_H491<=Vw;
XbG_H492<=Vw;
XbG_H493<=Vw;
XbG_H494<=Vw;
XbG_H495<=Vw;
XbG_H496<=Vw;
XbG_H497<=Vw;
XbG_H498<=Vw;
XbG_H499<=Vw;
XbG_H5<=Vw;
XbG_H50<=Vw;
XbG_H500<=Vw;
XbG_H501<=Vw;
XbG_H502<=Vw;
XbG_H503<=Vw;
XbG_H504<=Vw;
XbG_H505<=Vw;
XbG_H506<=Vw;
XbG_H507<=Vw;
XbG_H508<=Vw;
XbG_H509<=Vw;
XbG_H51<=Vw;
XbG_H510<=Vw;
XbG_H511<=Vw;
XbG_H512<=Vw;
XbG_H513<=Vw;
XbG_H514<=Vw;
XbG_H515<=Vw;
XbG_H516<=Vw;
XbG_H517<=Vw;
XbG_H518<=Vw;
XbG_H519<=Vw;
XbG_H52<=Vw;
XbG_H520<=Vw;
XbG_H521<=Vw;
XbG_H522<=Vw;
XbG_H523<=Vw;
XbG_H524<=Vw;
XbG_H525<=Vw;
XbG_H526<=Vw;
XbG_H527<=Vw;
XbG_H528<=Vw;
XbG_H529<=Vw;
XbG_H53<=Vw;
XbG_H530<=Vw;
XbG_H531<=Vw;
XbG_H532<=Vw;
XbG_H533<=Vw;
XbG_H534<=Vw;
XbG_H535<=Vw;
XbG_H536<=Vw;
XbG_H537<=Vw;
XbG_H538<=Vw;
XbG_H539<=Vw;
XbG_H54<=Vw;
XbG_H540<=Vw;
XbG_H541<=Vw;
XbG_H542<=Vw;
XbG_H543<=Vw;
XbG_H544<=Vw;
XbG_H545<=Vw;
XbG_H546<=Vw;
XbG_H547<=Vw;
XbG_H548<=Vw;
XbG_H549<=Vw;
XbG_H55<=Vw;
XbG_H550<=Vw;
XbG_H551<=Vw;
XbG_H552<=Vw;
XbG_H553<=Vw;
XbG_H554<=Vw;
XbG_H555<=Vw;
XbG_H556<=Vw;
XbG_H557<=Vw;
XbG_H558<=Vw;
XbG_H559<=Vw;
XbG_H56<=Vw;
XbG_H560<=Vw;
XbG_H561<=Vw;
XbG_H562<=Vw;
XbG_H563<=Vw;
XbG_H564<=Vw;
XbG_H565<=Vw;
XbG_H566<=Vw;
XbG_H567<=Vw;
XbG_H568<=Vw;
XbG_H569<=Vw;
XbG_H57<=Vw;
XbG_H570<=Vw;
XbG_H571<=Vw;
XbG_H572<=Vw;
XbG_H573<=Vw;
XbG_H574<=Vw;
XbG_H575<=Vw;
XbG_H576<=Vw;
XbG_H577<=Vw;
XbG_H578<=Vw;
XbG_H579<=Vw;
XbG_H58<=Vw;
XbG_H580<=Vw;
XbG_H581<=Vw;
XbG_H582<=Vw;
XbG_H583<=Vw;
XbG_H584<=Vw;
XbG_H585<=Vw;
XbG_H586<=Vw;
XbG_H587<=Vw;
XbG_H588<=Vw;
XbG_H589<=Vw;
XbG_H59<=Vw;
XbG_H590<=Vw;
XbG_H591<=Vw;
XbG_H592<=Vw;
XbG_H593<=Vw;
XbG_H594<=Vw;
XbG_H595<=Vw;
XbG_H596<=Vw;
XbG_H597<=Vw;
XbG_H598<=Vw;
XbG_H599<=Vw;
XbG_H6<=Vw;
XbG_H60<=Vw;
XbG_H600<=Vw;
XbG_H601<=Vw;
XbG_H602<=Vw;
XbG_H603<=Vw;
XbG_H604<=Vw;
XbG_H605<=Vw;
XbG_H606<=Vw;
XbG_H607<=Vw;
XbG_H608<=Vw;
XbG_H609<=Vw;
XbG_H61<=Vw;
XbG_H610<=Vw;
XbG_H611<=Vw;
XbG_H612<=Vw;
XbG_H613<=Vw;
XbG_H614<=Vw;
XbG_H615<=Vw;
XbG_H616<=Vw;
XbG_H617<=Vw;
XbG_H618<=Vw;
XbG_H619<=Vw;
XbG_H62<=Vw;
XbG_H620<=Vw;
XbG_H621<=Vw;
XbG_H622<=Vw;
XbG_H623<=Vw;
XbG_H624<=Vw;
XbG_H625<=Vw;
XbG_H626<=Vw;
XbG_H627<=Vw;
XbG_H628<=Vw;
XbG_H629<=Vw;
XbG_H63<=Vw;
XbG_H630<=Vw;
XbG_H631<=Vw;
XbG_H632<=Vw;
XbG_H633<=Vw;
XbG_H634<=Vw;
XbG_H635<=Vw;
XbG_H636<=Vw;
XbG_H637<=Vw;
XbG_H638<=Vw;
XbG_H639<=Vw;
XbG_H64<=Vw;
XbG_H640<=Vw;
XbG_H641<=Vw;
XbG_H642<=Vw;
XbG_H643<=Vw;
XbG_H644<=Vw;
XbG_H645<=Vw;
XbG_H646<=Vw;
XbG_H647<=Vw;
XbG_H648<=Vw;
XbG_H649<=Vw;
XbG_H65<=Vw;
XbG_H650<=Vw;
XbG_H651<=Vw;
XbG_H652<=Vw;
XbG_H653<=Vw;
XbG_H654<=Vw;
XbG_H655<=Vw;
XbG_H656<=Vw;
XbG_H657<=Vw;
XbG_H658<=Vw;
XbG_H659<=Vw;
XbG_H66<=Vw;
XbG_H660<=Vw;
XbG_H661<=Vw;
XbG_H662<=Vw;
XbG_H663<=Vw;
XbG_H664<=Vw;
XbG_H665<=Vw;
XbG_H666<=Vw;
XbG_H667<=Vw;
XbG_H668<=Vw;
XbG_H669<=Vw;
XbG_H67<=Vw;
XbG_H670<=Vw;
XbG_H671<=Vw;
XbG_H672<=Vw;
XbG_H673<=Vw;
XbG_H674<=Vw;
XbG_H675<=Vw;
XbG_H676<=Vw;
XbG_H677<=Vw;
XbG_H678<=Vw;
XbG_H679<=Vw;
XbG_H68<=Vw;
XbG_H680<=Vw;
XbG_H681<=Vw;
XbG_H682<=Vw;
XbG_H683<=Vw;
XbG_H684<=Vw;
XbG_H685<=Vw;
XbG_H686<=Vw;
XbG_H687<=Vw;
XbG_H688<=Vw;
XbG_H689<=Vw;
XbG_H69<=Vw;
XbG_H690<=Vw;
XbG_H691<=Vw;
XbG_H692<=Vw;
XbG_H693<=Vw;
XbG_H694<=Vw;
XbG_H695<=Vw;
XbG_H696<=Vw;
XbG_H697<=Vw;
XbG_H698<=Vw;
XbG_H699<=Vw;
XbG_H7<=Vw;
XbG_H70<=Vw;
XbG_H700<=Vw;
XbG_H701<=Vw;
XbG_H702<=Vw;
XbG_H703<=Vw;
XbG_H704<=Vw;
XbG_H705<=Vw;
XbG_H706<=Vw;
XbG_H707<=Vw;
XbG_H708<=Vw;
XbG_H709<=Vw;
XbG_H71<=Vw;
XbG_H710<=Vw;
XbG_H711<=Vw;
XbG_H712<=Vw;
XbG_H713<=Vw;
XbG_H714<=Vw;
XbG_H715<=Vw;
XbG_H716<=Vw;
XbG_H717<=Vw;
XbG_H718<=Vw;
XbG_H719<=Vw;
XbG_H72<=Vw;
XbG_H720<=Vw;
XbG_H721<=Vw;
XbG_H722<=Vr;
XbG_H723<=Vr;
XbG_H724<=Vr;
XbG_H725<=Vr;
XbG_H726<=Vr;
XbG_H727<=Vr;
XbG_H728<=Vr;
XbG_H729<=Vr;
XbG_H73<=Vw;
XbG_H730<=Vr;
XbG_H731<=Vr;
XbG_H732<=Vr;
XbG_H733<=Vr;
XbG_H734<=Vr;
XbG_H735<=Vr;
XbG_H74<=Vw;
XbG_H75<=Vw;
XbG_H76<=Vw;
XbG_H77<=Vw;
XbG_H78<=Vw;
XbG_H79<=Vw;
XbG_H8<=Vw;
XbG_H80<=Vw;
XbG_H81<=Vw;
XbG_H82<=Vw;
XbG_H83<=Vw;
XbG_H84<=Vw;
XbG_H85<=Vw;
XbG_H86<=Vw;
XbG_H87<=Vw;
XbG_H88<=Vw;
XbG_H89<=Vw;
XbG_H9<=Vw;
XbG_H90<=Vw;
XbG_H91<=Vw;
XbG_H92<=Vw;
XbG_H93<=Vw;
XbG_H94<=Vw;
XbG_H95<=Vw;
XbG_H96<=Vw;
XbG_H97<=Vw;
XbG_H98<=Vw;
XbG_H99<=Vw;
XbG_V0<=zero;
XbG_V1<=zero;
XbG_V10<=zero;
XbG_V100<=zero;
XbG_V101<=zero;
XbG_V102<=zero;
XbG_V103<=zero;
XbG_V104<=zero;
XbG_V105<=zero;
XbG_V106<=zero;
XbG_V107<=zero;
XbG_V108<=zero;
XbG_V109<=zero;
XbG_V11<=zero;
XbG_V110<=zero;
XbG_V111<=zero;
XbG_V112<=zero;
XbG_V113<=zero;
XbG_V114<=zero;
XbG_V115<=zero;
XbG_V116<=zero;
XbG_V117<=zero;
XbG_V118<=zero;
XbG_V119<=zero;
XbG_V12<=zero;
XbG_V120<=zero;
XbG_V121<=zero;
XbG_V122<=zero;
XbG_V123<=zero;
XbG_V124<=zero;
XbG_V125<=zero;
XbG_V126<=zero;
XbG_V127<=zero;
XbG_V128<=zero;
XbG_V129<=zero;
XbG_V13<=zero;
XbG_V130<=zero;
XbG_V131<=zero;
XbG_V132<=zero;
XbG_V133<=zero;
XbG_V134<=zero;
XbG_V135<=zero;
XbG_V136<=zero;
XbG_V137<=zero;
XbG_V138<=zero;
XbG_V139<=zero;
XbG_V14<=zero;
XbG_V140<=zero;
XbG_V141<=zero;
XbG_V142<=zero;
XbG_V143<=zero;
XbG_V144<=zero;
XbG_V145<=zero;
XbG_V146<=zero;
XbG_V147<=zero;
XbG_V148<=zero;
XbG_V149<=zero;
XbG_V15<=zero;
XbG_V150<=zero;
XbG_V151<=zero;
XbG_V152<=zero;
XbG_V153<=zero;
XbG_V154<=zero;
XbG_V155<=zero;
XbG_V156<=zero;
XbG_V157<=zero;
XbG_V158<=zero;
XbG_V159<=zero;
XbG_V16<=zero;
XbG_V160<=zero;
XbG_V161<=zero;
XbG_V162<=zero;
XbG_V163<=zero;
XbG_V164<=zero;
XbG_V165<=zero;
XbG_V166<=zero;
XbG_V167<=zero;
XbG_V168<=zero;
XbG_V169<=zero;
XbG_V17<=zero;
XbG_V170<=zero;
XbG_V171<=zero;
XbG_V172<=zero;
XbG_V173<=zero;
XbG_V174<=zero;
XbG_V175<=zero;
XbG_V176<=zero;
XbG_V177<=zero;
XbG_V178<=zero;
XbG_V179<=zero;
XbG_V18<=zero;
XbG_V180<=zero;
XbG_V181<=zero;
XbG_V182<=zero;
XbG_V183<=zero;
XbG_V184<=zero;
XbG_V185<=zero;
XbG_V186<=zero;
XbG_V187<=zero;
XbG_V188<=zero;
XbG_V189<=zero;
XbG_V19<=zero;
XbG_V2<=zero;
XbG_V20<=zero;
XbG_V21<=zero;
XbG_V22<=zero;
XbG_V23<=zero;
XbG_V24<=zero;
XbG_V25<=zero;
XbG_V26<=zero;
XbG_V27<=zero;
XbG_V28<=zero;
XbG_V29<=zero;
XbG_V3<=zero;
XbG_V30<=zero;
XbG_V31<=zero;
XbG_V32<=zero;
XbG_V33<=zero;
XbG_V34<=zero;
XbG_V35<=zero;
XbG_V36<=zero;
XbG_V37<=zero;
XbG_V38<=zero;
XbG_V39<=zero;
XbG_V4<=zero;
XbG_V40<=zero;
XbG_V41<=zero;
XbG_V42<=zero;
XbG_V43<=zero;
XbG_V44<=zero;
XbG_V45<=zero;
XbG_V46<=zero;
XbG_V47<=zero;
XbG_V48<=zero;
XbG_V49<=zero;
XbG_V5<=zero;
XbG_V50<=zero;
XbG_V51<=zero;
XbG_V52<=zero;
XbG_V53<=zero;
XbG_V54<=zero;
XbG_V55<=zero;
XbG_V56<=zero;
XbG_V57<=zero;
XbG_V58<=zero;
XbG_V59<=zero;
XbG_V6<=zero;
XbG_V60<=zero;
XbG_V61<=zero;
XbG_V62<=zero;
XbG_V63<=zero;
XbG_V64<=zero;
XbG_V65<=zero;
XbG_V66<=zero;
XbG_V67<=zero;
XbG_V68<=zero;
XbG_V69<=zero;
XbG_V7<=zero;
XbG_V70<=zero;
XbG_V71<=zero;
XbG_V72<=zero;
XbG_V73<=zero;
XbG_V74<=zero;
XbG_V75<=zero;
XbG_V76<=zero;
XbG_V77<=zero;
XbG_V78<=zero;
XbG_V79<=zero;
XbG_V8<=zero;
XbG_V80<=zero;
XbG_V81<=zero;
XbG_V82<=zero;
XbG_V83<=zero;
XbG_V84<=zero;
XbG_V85<=zero;
XbG_V86<=zero;
XbG_V87<=zero;
XbG_V88<=zero;
XbG_V89<=zero;
XbG_V9<=zero;
XbG_V90<=zero;
XbG_V91<=zero;
XbG_V92<=zero;
XbG_V93<=zero;
XbG_V94<=zero;
XbG_V95<=zero;
XbG_V96<=zero;
XbG_V97<=zero;
XbG_V98<=zero;
XbG_V99<=zero;

end if;

next_state<=B_RI;

when B_RI =>

XbG_H0<=zero;
XbG_H1<=Vr;
XbG_H2<=Vr;
XbG_H3<=Vr;
XbG_H4<=Vr;
XbG_H5<=Vr;
XbG_H6<=Vr;
XbG_H7<=Vr;
XbG_H8<=Vr;
XbG_H9<=Vr;
XbG_H10<=Vr;
XbG_H11<=Vr;
XbG_H12<=Vr;
XbG_H13<=Vr;
XbG_H14<=Vr;
XbG_H15<=Vr;
XbG_H16<=Vr;
XbG_H17<=Vr;
XbG_H18<=Vr;
XbG_H19<=Vr;
XbG_H20<=Vr;
XbG_H21<=Vr;
XbG_H22<=Vr;
XbG_H23<=Vr;
XbG_H24<=Vr;
XbG_H25<=Vr;
XbG_H26<=Vr;
XbG_H27<=Vr;
XbG_H28<=Vr;
XbG_H29<=Vr;
XbG_H30<=Vr;
XbG_H31<=Vr;
XbG_H32<=Vr;
XbG_H33<=Vr;
XbG_H34<=Vr;
XbG_H35<=Vr;
XbG_H36<=Vr;
XbG_H37<=Vr;
XbG_H38<=Vr;
XbG_H39<=Vr;
XbG_H40<=Vr;
XbG_H41<=Vr;
XbG_H42<=Vr;
XbG_H43<=Vr;
XbG_H44<=Vr;
XbG_H45<=Vr;
XbG_H46<=Vr;
XbG_H47<=Vr;
XbG_H48<=Vr;
XbG_H49<=Vr;
XbG_H50<=Vr;
XbG_H51<=Vr;
XbG_H52<=Vr;
XbG_H53<=Vr;
XbG_H54<=Vr;
XbG_H55<=Vr;
XbG_H56<=Vr;
XbG_H57<=Vr;
XbG_H58<=Vr;
XbG_H59<=Vr;
XbG_H60<=Vr;
XbG_H61<=Vr;
XbG_H62<=Vr;
XbG_H63<=Vr;
XbG_H64<=Vr;
XbG_H65<=Vr;
XbG_H66<=Vr;
XbG_H67<=Vr;
XbG_H68<=Vr;
XbG_H69<=Vr;
XbG_H70<=Vr;
XbG_H71<=Vr;
XbG_H72<=Vr;
XbG_H73<=Vr;
XbG_H74<=Vr;
XbG_H75<=Vr;
XbG_H76<=Vr;
XbG_H77<=Vr;
XbG_H78<=Vr;
XbG_H79<=Vr;
XbG_H80<=Vr;
XbG_H81<=Vr;
XbG_H82<=Vr;
XbG_H83<=Vr;
XbG_H84<=Vr;
XbG_H85<=Vr;
XbG_H86<=Vr;
XbG_H87<=Vr;
XbG_H88<=Vr;
XbG_H89<=Vr;
XbG_H90<=Vr;
XbG_H91<=Vr;
XbG_H92<=Vr;
XbG_H93<=Vr;
XbG_H94<=Vr;
XbG_H95<=Vr;
XbG_H96<=Vr;
XbG_H97<=Vr;
XbG_H98<=Vr;
XbG_H99<=Vr;
XbG_H100<=Vr;
XbG_H101<=Vr;
XbG_H102<=Vr;
XbG_H103<=Vr;
XbG_H104<=Vr;
XbG_H105<=Vr;
XbG_H106<=Vr;
XbG_H107<=Vr;
XbG_H108<=Vr;
XbG_H109<=Vr;
XbG_H110<=Vr;
XbG_H111<=Vr;
XbG_H112<=Vr;
XbG_H113<=Vr;
XbG_H114<=Vr;
XbG_H115<=Vr;
XbG_H116<=Vr;
XbG_H117<=Vr;
XbG_H118<=Vr;
XbG_H119<=Vr;
XbG_H120<=Vr;
XbG_H121<=Vr;
XbG_H122<=Vr;
XbG_H123<=Vr;
XbG_H124<=Vr;
XbG_H125<=Vr;
XbG_H126<=Vr;
XbG_H127<=Vr;
XbG_H128<=Vr;
XbG_H129<=Vr;
XbG_H130<=Vr;
XbG_H131<=Vr;
XbG_H132<=Vr;
XbG_H133<=Vr;
XbG_H134<=Vr;
XbG_H135<=Vr;
XbG_H136<=Vr;
XbG_H137<=Vr;
XbG_H138<=Vr;
XbG_H139<=Vr;
XbG_H140<=Vr;
XbG_H141<=Vr;
XbG_H142<=Vr;
XbG_H143<=Vr;
XbG_H144<=Vr;
XbG_H145<=Vr;
XbG_H146<=Vr;
XbG_H147<=Vr;
XbG_H148<=Vr;
XbG_H149<=Vr;
XbG_H150<=Vr;
XbG_H151<=Vr;
XbG_H152<=Vr;
XbG_H153<=Vr;
XbG_H154<=Vr;
XbG_H155<=Vr;
XbG_H156<=Vr;
XbG_H157<=Vr;
XbG_H158<=Vr;
XbG_H159<=Vr;
XbG_H160<=Vr;
XbG_H161<=Vr;
XbG_H162<=Vr;
XbG_H163<=Vr;
XbG_H164<=Vr;
XbG_H165<=Vr;
XbG_H166<=Vr;
XbG_H167<=Vr;
XbG_H168<=Vr;
XbG_H169<=Vr;
XbG_H170<=Vr;
XbG_H171<=Vr;
XbG_H172<=Vr;
XbG_H173<=Vr;
XbG_H174<=Vr;
XbG_H175<=Vr;
XbG_H176<=Vr;
XbG_H177<=Vr;
XbG_H178<=Vr;
XbG_H179<=Vr;
XbG_H180<=Vr;
XbG_H181<=Vr;
XbG_H182<=Vr;
XbG_H183<=Vr;
XbG_H184<=Vr;
XbG_H185<=Vr;
XbG_H186<=Vr;
XbG_H187<=Vr;
XbG_H188<=Vr;
XbG_H189<=Vr;
XbG_H190<=Vr;
XbG_H191<=Vr;
XbG_H192<=Vr;
XbG_H193<=Vr;
XbG_H194<=Vr;
XbG_H195<=Vr;
XbG_H196<=Vr;
XbG_H197<=Vr;
XbG_H198<=Vr;
XbG_H199<=Vr;
XbG_H200<=Vr;
XbG_H201<=Vr;
XbG_H202<=Vr;
XbG_H203<=Vr;
XbG_H204<=Vr;
XbG_H205<=Vr;
XbG_H206<=Vr;
XbG_H207<=Vr;
XbG_H208<=Vr;
XbG_H209<=Vr;
XbG_H210<=Vr;
XbG_H211<=Vr;
XbG_H212<=Vr;
XbG_H213<=Vr;
XbG_H214<=Vr;
XbG_H215<=Vr;
XbG_H216<=Vr;
XbG_H217<=Vr;
XbG_H218<=Vr;
XbG_H219<=Vr;
XbG_H220<=Vr;
XbG_H221<=Vr;
XbG_H222<=Vr;
XbG_H223<=Vr;
XbG_H224<=Vr;
XbG_H225<=Vr;
XbG_H226<=Vr;
XbG_H227<=Vr;
XbG_H228<=Vr;
XbG_H229<=Vr;
XbG_H230<=Vr;
XbG_H231<=Vr;
XbG_H232<=Vr;
XbG_H233<=Vr;
XbG_H234<=Vr;
XbG_H235<=Vr;
XbG_H236<=Vr;
XbG_H237<=Vr;
XbG_H238<=Vr;
XbG_H239<=Vr;
XbG_H240<=Vr;
XbG_H241<=Vr;
XbG_H242<=Vr;
XbG_H243<=Vr;
XbG_H244<=Vr;
XbG_H245<=Vr;
XbG_H246<=Vr;
XbG_H247<=Vr;
XbG_H248<=Vr;
XbG_H249<=Vr;
XbG_H250<=Vr;
XbG_H251<=Vr;
XbG_H252<=Vr;
XbG_H253<=Vr;
XbG_H254<=Vr;
XbG_H255<=Vr;
XbG_H256<=Vr;
XbG_H257<=Vr;
XbG_H258<=Vr;
XbG_H259<=Vr;
XbG_H260<=Vr;
XbG_H261<=Vr;
XbG_H262<=Vr;
XbG_H263<=Vr;
XbG_H264<=Vr;
XbG_H265<=Vr;
XbG_H266<=Vr;
XbG_H267<=Vr;
XbG_H268<=Vr;
XbG_H269<=Vr;
XbG_H270<=Vr;
XbG_H271<=Vr;
XbG_H272<=Vr;
XbG_H273<=Vr;
XbG_H274<=Vr;
XbG_H275<=Vr;
XbG_H276<=Vr;
XbG_H277<=Vr;
XbG_H278<=Vr;
XbG_H279<=Vr;
XbG_H280<=Vr;
XbG_H281<=Vr;
XbG_H282<=Vr;
XbG_H283<=Vr;
XbG_H284<=Vr;
XbG_H285<=Vr;
XbG_H286<=Vr;
XbG_H287<=Vr;
XbG_H288<=Vr;
XbG_H289<=Vr;
XbG_H290<=Vr;
XbG_H291<=Vr;
XbG_H292<=Vr;
XbG_H293<=Vr;
XbG_H294<=Vr;
XbG_H295<=Vr;
XbG_H296<=Vr;
XbG_H297<=Vr;
XbG_H298<=Vr;
XbG_H299<=Vr;
XbG_H300<=Vr;
XbG_H301<=Vr;
XbG_H302<=Vr;
XbG_H303<=Vr;
XbG_H304<=Vr;
XbG_H305<=Vr;
XbG_H306<=Vr;
XbG_H307<=Vr;
XbG_H308<=Vr;
XbG_H309<=Vr;
XbG_H310<=Vr;
XbG_H311<=Vr;
XbG_H312<=Vr;
XbG_H313<=Vr;
XbG_H314<=Vr;
XbG_H315<=Vr;
XbG_H316<=Vr;
XbG_H317<=Vr;
XbG_H318<=Vr;
XbG_H319<=Vr;
XbG_H320<=Vr;
XbG_H321<=Vr;
XbG_H322<=Vr;
XbG_H323<=Vr;
XbG_H324<=Vr;
XbG_H325<=Vr;
XbG_H326<=Vr;
XbG_H327<=Vr;
XbG_H328<=Vr;
XbG_H329<=Vr;
XbG_H330<=Vr;
XbG_H331<=Vr;
XbG_H332<=Vr;
XbG_H333<=Vr;
XbG_H334<=Vr;
XbG_H335<=Vr;
XbG_H336<=Vr;
XbG_H337<=Vr;
XbG_H338<=Vr;
XbG_H339<=Vr;
XbG_H340<=Vr;
XbG_H341<=Vr;
XbG_H342<=Vr;
XbG_H343<=Vr;
XbG_H344<=Vr;
XbG_H345<=Vr;
XbG_H346<=Vr;
XbG_H347<=Vr;
XbG_H348<=Vr;
XbG_H349<=Vr;
XbG_H350<=Vr;
XbG_H351<=Vr;
XbG_H352<=Vr;
XbG_H353<=Vr;
XbG_H354<=Vr;
XbG_H355<=Vr;
XbG_H356<=Vr;
XbG_H357<=Vr;
XbG_H358<=Vr;
XbG_H359<=Vr;
XbG_H360<=Vr;
XbG_H361<=Vr;
XbG_H362<=Vr;
XbG_H363<=Vr;
XbG_H364<=Vr;
XbG_H365<=Vr;
XbG_H366<=Vr;
XbG_H367<=Vr;
XbG_H368<=Vr;
XbG_H369<=Vr;
XbG_H370<=Vr;
XbG_H371<=Vr;
XbG_H372<=Vr;
XbG_H373<=Vr;
XbG_H374<=Vr;
XbG_H375<=Vr;
XbG_H376<=Vr;
XbG_H377<=Vr;
XbG_H378<=Vr;
XbG_H379<=Vr;
XbG_H380<=Vr;
XbG_H381<=Vr;
XbG_H382<=Vr;
XbG_H383<=Vr;
XbG_H384<=Vr;
XbG_H385<=Vr;
XbG_H386<=Vr;
XbG_H387<=Vr;
XbG_H388<=Vr;
XbG_H389<=Vr;
XbG_H390<=Vr;
XbG_H391<=Vr;
XbG_H392<=Vr;
XbG_H393<=Vr;
XbG_H394<=Vr;
XbG_H395<=Vr;
XbG_H396<=Vr;
XbG_H397<=Vr;
XbG_H398<=Vr;
XbG_H399<=Vr;
XbG_H400<=Vr;
XbG_H401<=Vr;
XbG_H402<=Vr;
XbG_H403<=Vr;
XbG_H404<=Vr;
XbG_H405<=Vr;
XbG_H406<=Vr;
XbG_H407<=Vr;
XbG_H408<=Vr;
XbG_H409<=Vr;
XbG_H410<=Vr;
XbG_H411<=Vr;
XbG_H412<=Vr;
XbG_H413<=Vr;
XbG_H414<=Vr;
XbG_H415<=Vr;
XbG_H416<=Vr;
XbG_H417<=Vr;
XbG_H418<=Vr;
XbG_H419<=Vr;
XbG_H420<=Vr;
XbG_H421<=Vr;
XbG_H422<=Vr;
XbG_H423<=Vr;
XbG_H424<=Vr;
XbG_H425<=Vr;
XbG_H426<=Vr;
XbG_H427<=Vr;
XbG_H428<=Vr;
XbG_H429<=Vr;
XbG_H430<=Vr;
XbG_H431<=Vr;
XbG_H432<=Vr;
XbG_H433<=Vr;
XbG_H434<=Vr;
XbG_H435<=Vr;
XbG_H436<=Vr;
XbG_H437<=Vr;
XbG_H438<=Vr;
XbG_H439<=Vr;
XbG_H440<=Vr;
XbG_H441<=Vr;
XbG_H442<=Vr;
XbG_H443<=Vr;
XbG_H444<=Vr;
XbG_H445<=Vr;
XbG_H446<=Vr;
XbG_H447<=Vr;
XbG_H448<=Vr;
XbG_H449<=Vr;
XbG_H450<=Vr;
XbG_H451<=Vr;
XbG_H452<=Vr;
XbG_H453<=Vr;
XbG_H454<=Vr;
XbG_H455<=Vr;
XbG_H456<=Vr;
XbG_H457<=Vr;
XbG_H458<=Vr;
XbG_H459<=Vr;
XbG_H460<=Vr;
XbG_H461<=Vr;
XbG_H462<=Vr;
XbG_H463<=Vr;
XbG_H464<=Vr;
XbG_H465<=Vr;
XbG_H466<=Vr;
XbG_H467<=Vr;
XbG_H468<=Vr;
XbG_H469<=Vr;
XbG_H470<=Vr;
XbG_H471<=Vr;
XbG_H472<=Vr;
XbG_H473<=Vr;
XbG_H474<=Vr;
XbG_H475<=Vr;
XbG_H476<=Vr;
XbG_H477<=Vr;
XbG_H478<=Vr;
XbG_H479<=Vr;
XbG_H480<=Vr;
XbG_H481<=Vr;
XbG_H482<=Vr;
XbG_H483<=Vr;
XbG_H484<=Vr;
XbG_H485<=Vr;
XbG_H486<=Vr;
XbG_H487<=Vr;
XbG_H488<=Vr;
XbG_H489<=Vr;
XbG_H490<=Vr;
XbG_H491<=Vr;
XbG_H492<=Vr;
XbG_H493<=Vr;
XbG_H494<=Vr;
XbG_H495<=Vr;
XbG_H496<=Vr;
XbG_H497<=Vr;
XbG_H498<=Vr;
XbG_H499<=Vr;
XbG_H500<=Vr;
XbG_H501<=Vr;
XbG_H502<=Vr;
XbG_H503<=Vr;
XbG_H504<=Vr;
XbG_H505<=Vr;
XbG_H506<=Vr;
XbG_H507<=Vr;
XbG_H508<=Vr;
XbG_H509<=Vr;
XbG_H510<=Vr;
XbG_H511<=Vr;
XbG_H512<=Vr;
XbG_H513<=Vr;
XbG_H514<=Vr;
XbG_H515<=Vr;
XbG_H516<=Vr;
XbG_H517<=Vr;
XbG_H518<=Vr;
XbG_H519<=Vr;
XbG_H520<=Vr;
XbG_H521<=Vr;
XbG_H522<=Vr;
XbG_H523<=Vr;
XbG_H524<=Vr;
XbG_H525<=Vr;
XbG_H526<=Vr;
XbG_H527<=Vr;
XbG_H528<=Vr;
XbG_H529<=Vr;
XbG_H530<=Vr;
XbG_H531<=Vr;
XbG_H532<=Vr;
XbG_H533<=Vr;
XbG_H534<=Vr;
XbG_H535<=Vr;
XbG_H536<=Vr;
XbG_H537<=Vr;
XbG_H538<=Vr;
XbG_H539<=Vr;
XbG_H540<=Vr;
XbG_H541<=Vr;
XbG_H542<=Vr;
XbG_H543<=Vr;
XbG_H544<=Vr;
XbG_H545<=Vr;
XbG_H546<=Vr;
XbG_H547<=Vr;
XbG_H548<=Vr;
XbG_H549<=Vr;
XbG_H550<=Vr;
XbG_H551<=Vr;
XbG_H552<=Vr;
XbG_H553<=Vr;
XbG_H554<=Vr;
XbG_H555<=Vr;
XbG_H556<=Vr;
XbG_H557<=Vr;
XbG_H558<=Vr;
XbG_H559<=Vr;
XbG_H560<=Vr;
XbG_H561<=Vr;
XbG_H562<=Vr;
XbG_H563<=Vr;
XbG_H564<=Vr;
XbG_H565<=Vr;
XbG_H566<=Vr;
XbG_H567<=Vr;
XbG_H568<=Vr;
XbG_H569<=Vr;
XbG_H570<=Vr;
XbG_H571<=Vr;
XbG_H572<=Vr;
XbG_H573<=Vr;
XbG_H574<=Vr;
XbG_H575<=Vr;
XbG_H576<=Vr;
XbG_H577<=Vr;
XbG_H578<=Vr;
XbG_H579<=Vr;
XbG_H580<=Vr;
XbG_H581<=Vr;
XbG_H582<=Vr;
XbG_H583<=Vr;
XbG_H584<=Vr;
XbG_H585<=Vr;
XbG_H586<=Vr;
XbG_H587<=Vr;
XbG_H588<=Vr;
XbG_H589<=Vr;
XbG_H590<=Vr;
XbG_H591<=Vr;
XbG_H592<=Vr;
XbG_H593<=Vr;
XbG_H594<=Vr;
XbG_H595<=Vr;
XbG_H596<=Vr;
XbG_H597<=Vr;
XbG_H598<=Vr;
XbG_H599<=Vr;
XbG_H600<=Vr;
XbG_H601<=Vr;
XbG_H602<=Vr;
XbG_H603<=Vr;
XbG_H604<=Vr;
XbG_H605<=Vr;
XbG_H606<=Vr;
XbG_H607<=Vr;
XbG_H608<=Vr;
XbG_H609<=Vr;
XbG_H610<=Vr;
XbG_H611<=Vr;
XbG_H612<=Vr;
XbG_H613<=Vr;
XbG_H614<=Vr;
XbG_H615<=Vr;
XbG_H616<=Vr;
XbG_H617<=Vr;
XbG_H618<=Vr;
XbG_H619<=Vr;
XbG_H620<=Vr;
XbG_H621<=Vr;
XbG_H622<=Vr;
XbG_H623<=Vr;
XbG_H624<=Vr;
XbG_H625<=Vr;
XbG_H626<=Vr;
XbG_H627<=Vr;
XbG_H628<=Vr;
XbG_H629<=Vr;
XbG_H630<=Vr;
XbG_H631<=Vr;
XbG_H632<=Vr;
XbG_H633<=Vr;
XbG_H634<=Vr;
XbG_H635<=Vr;
XbG_H636<=Vr;
XbG_H637<=Vr;
XbG_H638<=Vr;
XbG_H639<=Vr;
XbG_H640<=Vr;
XbG_H641<=Vr;
XbG_H642<=Vr;
XbG_H643<=Vr;
XbG_H644<=Vr;
XbG_H645<=Vr;
XbG_H646<=Vr;
XbG_H647<=Vr;
XbG_H648<=Vr;
XbG_H649<=Vr;
XbG_H650<=Vr;
XbG_H651<=Vr;
XbG_H652<=Vr;
XbG_H653<=Vr;
XbG_H654<=Vr;
XbG_H655<=Vr;
XbG_H656<=Vr;
XbG_H657<=Vr;
XbG_H658<=Vr;
XbG_H659<=Vr;
XbG_H660<=Vr;
XbG_H661<=Vr;
XbG_H662<=Vr;
XbG_H663<=Vr;
XbG_H664<=Vr;
XbG_H665<=Vr;
XbG_H666<=Vr;
XbG_H667<=Vr;
XbG_H668<=Vr;
XbG_H669<=Vr;
XbG_H670<=Vr;
XbG_H671<=Vr;
XbG_H672<=Vr;
XbG_H673<=Vr;
XbG_H674<=Vr;
XbG_H675<=Vr;
XbG_H676<=Vr;
XbG_H677<=Vr;
XbG_H678<=Vr;
XbG_H679<=Vr;
XbG_H680<=Vr;
XbG_H681<=Vr;
XbG_H682<=Vr;
XbG_H683<=Vr;
XbG_H684<=Vr;
XbG_H685<=Vr;
XbG_H686<=Vr;
XbG_H687<=Vr;
XbG_H688<=Vr;
XbG_H689<=Vr;
XbG_H690<=Vr;
XbG_H691<=Vr;
XbG_H692<=Vr;
XbG_H693<=Vr;
XbG_H694<=Vr;
XbG_H695<=Vr;
XbG_H696<=Vr;
XbG_H697<=Vr;
XbG_H698<=Vr;
XbG_H699<=Vr;
XbG_H700<=Vr;
XbG_H701<=Vr;
XbG_H702<=Vr;
XbG_H703<=Vr;
XbG_H704<=Vr;
XbG_H705<=Vr;
XbG_H706<=Vr;
XbG_H707<=Vr;
XbG_H708<=Vr;
XbG_H709<=Vr;
XbG_H710<=Vr;
XbG_H711<=Vr;
XbG_H712<=Vr;
XbG_H713<=Vr;
XbG_H714<=Vr;
XbG_H715<=Vr;
XbG_H716<=Vr;
XbG_H717<=Vr;
XbG_H718<=Vr;
XbG_H719<=Vr;
XbG_H720<=Vr;
XbG_H721<=Vr;

if pi26='1' then XbG_V0<=Vw_neg; else XbG_V0<=Vw; end if;

if pi26='0' then XbG_V1<=Vw_neg; else XbG_V1<=Vw; end if;

if pi15='1' then XbG_V2<=Vw_neg; else XbG_V2<=Vw; end if;

if pi15='0' then XbG_V3<=Vw_neg; else XbG_V3<=Vw; end if;

if pi00='1' then XbG_V18<=Vw_neg; else XbG_V18<=Vw; end if;

if pi00='0' then XbG_V19<=Vw_neg; else XbG_V19<=Vw; end if;

if pi06='1' then XbG_V20<=Vw_neg; else XbG_V20<=Vw; end if;

if pi06='0' then XbG_V21<=Vw_neg; else XbG_V21<=Vw; end if;

if pi03='1' then XbG_V22<=Vw_neg; else XbG_V22<=Vw; end if;

if pi03='0' then XbG_V23<=Vw_neg; else XbG_V23<=Vw; end if;

if pi07='1' then XbG_V24<=Vw_neg; else XbG_V24<=Vw; end if;

if pi07='0' then XbG_V25<=Vw_neg; else XbG_V25<=Vw; end if;

if pi08='1' then XbG_V26<=Vw_neg; else XbG_V26<=Vw; end if;

if pi08='0' then XbG_V27<=Vw_neg; else XbG_V27<=Vw; end if;

if pi09='1' then XbG_V28<=Vw_neg; else XbG_V28<=Vw; end if;

if pi09='0' then XbG_V29<=Vw_neg; else XbG_V29<=Vw; end if;

if pi10='1' then XbG_V30<=Vw_neg; else XbG_V30<=Vw; end if;

if pi10='0' then XbG_V31<=Vw_neg; else XbG_V31<=Vw; end if;

if pi02='1' then XbG_V32<=Vw_neg; else XbG_V32<=Vw; end if;

if pi02='0' then XbG_V33<=Vw_neg; else XbG_V33<=Vw; end if;

if pi17='1' then XbG_V34<=Vw_neg; else XbG_V34<=Vw; end if;

if pi17='0' then XbG_V35<=Vw_neg; else XbG_V35<=Vw; end if;

if pi01='1' then XbG_V36<=Vw_neg; else XbG_V36<=Vw; end if;

if pi01='0' then XbG_V37<=Vw_neg; else XbG_V37<=Vw; end if;

if pi11='1' then XbG_V38<=Vw_neg; else XbG_V38<=Vw; end if;

if pi11='0' then XbG_V39<=Vw_neg; else XbG_V39<=Vw; end if;

if pi12='1' then XbG_V40<=Vw_neg; else XbG_V40<=Vw; end if;

if pi12='0' then XbG_V41<=Vw_neg; else XbG_V41<=Vw; end if;

if pi13='1' then XbG_V42<=Vw_neg; else XbG_V42<=Vw; end if;

if pi13='0' then XbG_V43<=Vw_neg; else XbG_V43<=Vw; end if;

if pi14='1' then XbG_V44<=Vw_neg; else XbG_V44<=Vw; end if;

if pi14='0' then XbG_V45<=Vw_neg; else XbG_V45<=Vw; end if;

if pi04='1' then XbG_V46<=Vw_neg; else XbG_V46<=Vw; end if;

if pi04='0' then XbG_V47<=Vw_neg; else XbG_V47<=Vw; end if;

if pi16='1' then XbG_V48<=Vw_neg; else XbG_V48<=Vw; end if;

if pi16='0' then XbG_V49<=Vw_neg; else XbG_V49<=Vw; end if;

if pi05='1' then XbG_V50<=Vw_neg; else XbG_V50<=Vw; end if;

if pi05='0' then XbG_V51<=Vw_neg; else XbG_V51<=Vw; end if;

if pi18='1' then XbG_V52<=Vw_neg; else XbG_V52<=Vw; end if;

if pi18='0' then XbG_V53<=Vw_neg; else XbG_V53<=Vw; end if;

if pi19='1' then XbG_V54<=Vw_neg; else XbG_V54<=Vw; end if;

if pi19='0' then XbG_V55<=Vw_neg; else XbG_V55<=Vw; end if;

if pi20='1' then XbG_V56<=Vw_neg; else XbG_V56<=Vw; end if;

if pi20='0' then XbG_V57<=Vw_neg; else XbG_V57<=Vw; end if;

if pi21='1' then XbG_V58<=Vw_neg; else XbG_V58<=Vw; end if;

if pi21='0' then XbG_V59<=Vw_neg; else XbG_V59<=Vw; end if;

if pi22='1' then XbG_V60<=Vw_neg; else XbG_V60<=Vw; end if;

if pi22='0' then XbG_V61<=Vw_neg; else XbG_V61<=Vw; end if;

if pi23='1' then XbG_V62<=Vw_neg; else XbG_V62<=Vw; end if;

if pi23='0' then XbG_V63<=Vw_neg; else XbG_V63<=Vw; end if;

if pi24='1' then XbG_V64<=Vw_neg; else XbG_V64<=Vw; end if;

if pi24='0' then XbG_V65<=Vw_neg; else XbG_V65<=Vw; end if;

if pi25='1' then XbG_V66<=Vw_neg; else XbG_V66<=Vw; end if;

if pi25='0' then XbG_V67<=Vw_neg; else XbG_V67<=Vw; end if;

XbG_V68<=Vr;
XbG_V69<=Vr;
XbG_V70<=Vr;
XbG_V71<=Vr;
XbG_V72<=Vr;
XbG_V73<=Vr;
XbG_V74<=Vr;
XbG_V75<=Vr;
XbG_V76<=Vr;
XbG_V77<=Vr;
XbG_V78<=Vr;
XbG_V79<=Vr;
XbG_V80<=Vr;
XbG_V81<=Vr;
XbG_V82<=Vr;
XbG_V83<=Vr;
XbG_V84<=Vr;
XbG_V85<=Vr;
XbG_V86<=Vr;
XbG_V87<=Vr;
XbG_V88<=Vr;
XbG_V89<=Vr;
XbG_V90<=Vr;
XbG_V91<=Vr;
XbG_V92<=Vr;
XbG_V93<=Vr;
XbG_V94<=Vr;
XbG_V95<=Vr;
XbG_V96<=Vr;
XbG_V97<=Vr;
XbG_V98<=Vr;
XbG_V99<=Vr;
XbG_V100<=Vr;
XbG_V101<=Vr;
XbG_V102<=Vr;
XbG_V103<=Vr;
XbG_V104<=Vr;
XbG_V105<=Vr;
XbG_V106<=Vr;
XbG_V107<=Vr;
XbG_V108<=Vr;
XbG_V109<=Vr;
XbG_V110<=Vr;
XbG_V111<=Vr;
XbG_V112<=Vr;
XbG_V113<=Vr;
XbG_V114<=Vr;
XbG_V115<=Vr;
XbG_V116<=Vr;
XbG_V117<=Vr;
XbG_V118<=Vr;
XbG_V119<=Vr;
XbG_V120<=Vr;
XbG_V121<=Vr;
XbG_V122<=Vr;
XbG_V123<=Vr;
XbG_V124<=Vr;
XbG_V125<=Vr;
XbG_V126<=Vr;
XbG_V127<=Vr;
XbG_V128<=Vr;
XbG_V129<=Vr;
XbG_V130<=Vr;
XbG_V131<=Vr;
XbG_V132<=Vr;
XbG_V133<=Vr;
XbG_V134<=Vr;
XbG_V135<=Vr;
XbG_V136<=Vr;
XbG_V137<=Vr;
XbG_V138<=Vr;
XbG_V139<=Vr;
XbG_V140<=Vr;
XbG_V141<=Vr;
XbG_V142<=Vr;
XbG_V143<=Vr;
XbG_V144<=Vr;
XbG_V145<=Vr;
XbG_V146<=Vr;
XbG_V147<=Vr;
XbG_V148<=Vr;
XbG_V149<=Vr;
XbG_V150<=Vr;
XbG_V151<=Vr;
XbG_V152<=Vr;
XbG_V153<=Vr;
XbG_V154<=Vr;
XbG_V155<=Vr;
XbG_V156<=Vr;
XbG_V157<=Vr;
XbG_V158<=Vr;
XbG_V159<=Vr;
XbG_V160<=Vr;
XbG_V161<=Vr;
XbG_V162<=Vr;
XbG_V163<=Vr;
XbG_V164<=Vr;
XbG_V165<=Vr;
XbG_V166<=Vr;
XbG_V167<=Vr;
XbG_V168<=Vr;
XbG_V169<=Vr;
XbG_V170<=Vr;
XbG_V171<=Vr;
XbG_V172<=Vr;
XbG_V173<=Vr;
XbG_V174<=Vr;
XbG_V175<=Vr;
XbG_V176<=Vr;
XbG_V177<=Vr;
XbG_V178<=Vr;
XbG_V179<=Vr;
XbG_V180<=Vr;
XbG_V181<=Vr;
XbG_V182<=Vr;
XbG_V183<=Vr;
XbG_V184<=Vr;
XbG_V185<=Vr;
XbG_V186<=Vr;
XbG_V187<=Vr;
XbG_V188<=Vr;
XbG_V189<=Vr;

if feedback_enable = '0' then

if lo0='1' then XbG_V16<=Vw_neg; else XbG_V16<=Vw; end if;

if lo0='0' then XbG_V17<=Vw_neg; else XbG_V17<=Vw; end if;

if lo1='1' then XbG_V14<=Vw_neg; else XbG_V14<=Vw; end if;

if lo1='0' then XbG_V15<=Vw_neg; else XbG_V15<=Vw; end if;

if lo2='1' then XbG_V12<=Vw_neg; else XbG_V12<=Vw; end if;

if lo2='0' then XbG_V13<=Vw_neg; else XbG_V13<=Vw; end if;

if lo3='1' then XbG_V10<=Vw_neg; else XbG_V10<=Vw; end if;

if lo3='0' then XbG_V11<=Vw_neg; else XbG_V11<=Vw; end if;

if lo4='1' then XbG_V8<=Vw_neg; else XbG_V8<=Vw; end if;

if lo4='0' then XbG_V9<=Vw_neg; else XbG_V9<=Vw; end if;

if lo5='1' then XbG_V6<=Vw_neg; else XbG_V6<=Vw; end if;

if lo5='0' then XbG_V7<=Vw_neg; else XbG_V7<=Vw; end if;

if lo6='1' then XbG_V4<=Vw_neg; else XbG_V4<=Vw; end if;

if lo6='0' then XbG_V5<=Vw_neg; else XbG_V5<=Vw; end if;

XbG_H722<=zero;
XbG_H723<=zero;
XbG_H724<=zero;
XbG_H725<=zero;
XbG_H726<=zero;
XbG_H727<=zero;
XbG_H728<=zero;
XbG_H729<=zero;
XbG_H730<=zero;
XbG_H731<=zero;
XbG_H732<=zero;
XbG_H733<=zero;
XbG_H734<=zero;
XbG_H735<=zero;

else

XbG_V16<=Vw;
XbG_V17<=Vw;
XbG_V14<=Vw;
XbG_V15<=Vw;
XbG_V12<=Vw;
XbG_V13<=Vw;
XbG_V10<=Vw;
XbG_V11<=Vw;
XbG_V8<=Vw;
XbG_V9<=Vw;
XbG_V6<=Vw;
XbG_V7<=Vw;
XbG_V4<=Vw;
XbG_V5<=Vw;
XbG_H722<=zero, (others=>'Z') after 1 ps;
XbG_H723<=zero, (others=>'Z') after 1 ps;
XbG_H724<=zero, (others=>'Z') after 1 ps;
XbG_H725<=zero, (others=>'Z') after 1 ps;
XbG_H726<=zero, (others=>'Z') after 1 ps;
XbG_H727<=zero, (others=>'Z') after 1 ps;
XbG_H728<=zero, (others=>'Z') after 1 ps;
XbG_H729<=zero, (others=>'Z') after 1 ps;
XbG_H730<=zero, (others=>'Z') after 1 ps;
XbG_H731<=zero, (others=>'Z') after 1 ps;
XbG_H732<=zero, (others=>'Z') after 1 ps;
XbG_H733<=zero, (others=>'Z') after 1 ps;
XbG_H734<=zero, (others=>'Z') after 1 ps;
XbG_H735<=zero, (others=>'Z') after 1 ps;

end if;

next_state<=C_CFM;

when C_CFM =>

XbG_H0<=Vw;
XbG_H1<=zero;
XbG_H10<=zero;
XbG_H100<=zero;
XbG_H101<=zero;
XbG_H102<=zero;
XbG_H103<=zero;
XbG_H104<=zero;
XbG_H105<=zero;
XbG_H106<=zero;
XbG_H107<=zero;
XbG_H108<=zero;
XbG_H109<=zero;
XbG_H11<=zero;
XbG_H110<=zero;
XbG_H111<=zero;
XbG_H112<=zero;
XbG_H113<=zero;
XbG_H114<=zero;
XbG_H115<=zero;
XbG_H116<=zero;
XbG_H117<=zero;
XbG_H118<=zero;
XbG_H119<=zero;
XbG_H12<=zero;
XbG_H120<=zero;
XbG_H121<=zero;
XbG_H122<=zero;
XbG_H123<=zero;
XbG_H124<=zero;
XbG_H125<=zero;
XbG_H126<=zero;
XbG_H127<=zero;
XbG_H128<=zero;
XbG_H129<=zero;
XbG_H13<=zero;
XbG_H130<=zero;
XbG_H131<=zero;
XbG_H132<=zero;
XbG_H133<=zero;
XbG_H134<=zero;
XbG_H135<=zero;
XbG_H136<=zero;
XbG_H137<=zero;
XbG_H138<=zero;
XbG_H139<=zero;
XbG_H14<=zero;
XbG_H140<=zero;
XbG_H141<=zero;
XbG_H142<=zero;
XbG_H143<=zero;
XbG_H144<=zero;
XbG_H145<=zero;
XbG_H146<=zero;
XbG_H147<=zero;
XbG_H148<=zero;
XbG_H149<=zero;
XbG_H15<=zero;
XbG_H150<=zero;
XbG_H151<=zero;
XbG_H152<=zero;
XbG_H153<=zero;
XbG_H154<=zero;
XbG_H155<=zero;
XbG_H156<=zero;
XbG_H157<=zero;
XbG_H158<=zero;
XbG_H159<=zero;
XbG_H16<=zero;
XbG_H160<=zero;
XbG_H161<=zero;
XbG_H162<=zero;
XbG_H163<=zero;
XbG_H164<=zero;
XbG_H165<=zero;
XbG_H166<=zero;
XbG_H167<=zero;
XbG_H168<=zero;
XbG_H169<=zero;
XbG_H17<=zero;
XbG_H170<=zero;
XbG_H171<=zero;
XbG_H172<=zero;
XbG_H173<=zero;
XbG_H174<=zero;
XbG_H175<=zero;
XbG_H176<=zero;
XbG_H177<=zero;
XbG_H178<=zero;
XbG_H179<=zero;
XbG_H18<=zero;
XbG_H180<=zero;
XbG_H181<=zero;
XbG_H182<=zero;
XbG_H183<=zero;
XbG_H184<=zero;
XbG_H185<=zero;
XbG_H186<=zero;
XbG_H187<=zero;
XbG_H188<=zero;
XbG_H189<=zero;
XbG_H19<=zero;
XbG_H190<=zero;
XbG_H191<=zero;
XbG_H192<=zero;
XbG_H193<=zero;
XbG_H194<=zero;
XbG_H195<=zero;
XbG_H196<=zero;
XbG_H197<=zero;
XbG_H198<=zero;
XbG_H199<=zero;
XbG_H2<=zero;
XbG_H20<=zero;
XbG_H200<=zero;
XbG_H201<=zero;
XbG_H202<=zero;
XbG_H203<=zero;
XbG_H204<=zero;
XbG_H205<=zero;
XbG_H206<=zero;
XbG_H207<=zero;
XbG_H208<=zero;
XbG_H209<=zero;
XbG_H21<=zero;
XbG_H210<=zero;
XbG_H211<=zero;
XbG_H212<=zero;
XbG_H213<=zero;
XbG_H214<=zero;
XbG_H215<=zero;
XbG_H216<=zero;
XbG_H217<=zero;
XbG_H218<=zero;
XbG_H219<=zero;
XbG_H22<=zero;
XbG_H220<=zero;
XbG_H221<=zero;
XbG_H222<=zero;
XbG_H223<=zero;
XbG_H224<=zero;
XbG_H225<=zero;
XbG_H226<=zero;
XbG_H227<=zero;
XbG_H228<=zero;
XbG_H229<=zero;
XbG_H23<=zero;
XbG_H230<=zero;
XbG_H231<=zero;
XbG_H232<=zero;
XbG_H233<=zero;
XbG_H234<=zero;
XbG_H235<=zero;
XbG_H236<=zero;
XbG_H237<=zero;
XbG_H238<=zero;
XbG_H239<=zero;
XbG_H24<=zero;
XbG_H240<=zero;
XbG_H241<=zero;
XbG_H242<=zero;
XbG_H243<=zero;
XbG_H244<=zero;
XbG_H245<=zero;
XbG_H246<=zero;
XbG_H247<=zero;
XbG_H248<=zero;
XbG_H249<=zero;
XbG_H25<=zero;
XbG_H250<=zero;
XbG_H251<=zero;
XbG_H252<=zero;
XbG_H253<=zero;
XbG_H254<=zero;
XbG_H255<=zero;
XbG_H256<=zero;
XbG_H257<=zero;
XbG_H258<=zero;
XbG_H259<=zero;
XbG_H26<=zero;
XbG_H260<=zero;
XbG_H261<=zero;
XbG_H262<=zero;
XbG_H263<=zero;
XbG_H264<=zero;
XbG_H265<=zero;
XbG_H266<=zero;
XbG_H267<=zero;
XbG_H268<=zero;
XbG_H269<=zero;
XbG_H27<=zero;
XbG_H270<=zero;
XbG_H271<=zero;
XbG_H272<=zero;
XbG_H273<=zero;
XbG_H274<=zero;
XbG_H275<=zero;
XbG_H276<=zero;
XbG_H277<=zero;
XbG_H278<=zero;
XbG_H279<=zero;
XbG_H28<=zero;
XbG_H280<=zero;
XbG_H281<=zero;
XbG_H282<=zero;
XbG_H283<=zero;
XbG_H284<=zero;
XbG_H285<=zero;
XbG_H286<=zero;
XbG_H287<=zero;
XbG_H288<=zero;
XbG_H289<=zero;
XbG_H29<=zero;
XbG_H290<=zero;
XbG_H291<=zero;
XbG_H292<=zero;
XbG_H293<=zero;
XbG_H294<=zero;
XbG_H295<=zero;
XbG_H296<=zero;
XbG_H297<=zero;
XbG_H298<=zero;
XbG_H299<=zero;
XbG_H3<=zero;
XbG_H30<=zero;
XbG_H300<=zero;
XbG_H301<=zero;
XbG_H302<=zero;
XbG_H303<=zero;
XbG_H304<=zero;
XbG_H305<=zero;
XbG_H306<=zero;
XbG_H307<=zero;
XbG_H308<=zero;
XbG_H309<=zero;
XbG_H31<=zero;
XbG_H310<=zero;
XbG_H311<=zero;
XbG_H312<=zero;
XbG_H313<=zero;
XbG_H314<=zero;
XbG_H315<=zero;
XbG_H316<=zero;
XbG_H317<=zero;
XbG_H318<=zero;
XbG_H319<=zero;
XbG_H32<=zero;
XbG_H320<=zero;
XbG_H321<=zero;
XbG_H322<=zero;
XbG_H323<=zero;
XbG_H324<=zero;
XbG_H325<=zero;
XbG_H326<=zero;
XbG_H327<=zero;
XbG_H328<=zero;
XbG_H329<=zero;
XbG_H33<=zero;
XbG_H330<=zero;
XbG_H331<=zero;
XbG_H332<=zero;
XbG_H333<=zero;
XbG_H334<=zero;
XbG_H335<=zero;
XbG_H336<=zero;
XbG_H337<=zero;
XbG_H338<=zero;
XbG_H339<=zero;
XbG_H34<=zero;
XbG_H340<=zero;
XbG_H341<=zero;
XbG_H342<=zero;
XbG_H343<=zero;
XbG_H344<=zero;
XbG_H345<=zero;
XbG_H346<=zero;
XbG_H347<=zero;
XbG_H348<=zero;
XbG_H349<=zero;
XbG_H35<=zero;
XbG_H350<=zero;
XbG_H351<=zero;
XbG_H352<=zero;
XbG_H353<=zero;
XbG_H354<=zero;
XbG_H355<=zero;
XbG_H356<=zero;
XbG_H357<=zero;
XbG_H358<=zero;
XbG_H359<=zero;
XbG_H36<=zero;
XbG_H360<=zero;
XbG_H361<=zero;
XbG_H362<=zero;
XbG_H363<=zero;
XbG_H364<=zero;
XbG_H365<=zero;
XbG_H366<=zero;
XbG_H367<=zero;
XbG_H368<=zero;
XbG_H369<=zero;
XbG_H37<=zero;
XbG_H370<=zero;
XbG_H371<=zero;
XbG_H372<=zero;
XbG_H373<=zero;
XbG_H374<=zero;
XbG_H375<=zero;
XbG_H376<=zero;
XbG_H377<=zero;
XbG_H378<=zero;
XbG_H379<=zero;
XbG_H38<=zero;
XbG_H380<=zero;
XbG_H381<=zero;
XbG_H382<=zero;
XbG_H383<=zero;
XbG_H384<=zero;
XbG_H385<=zero;
XbG_H386<=zero;
XbG_H387<=zero;
XbG_H388<=zero;
XbG_H389<=zero;
XbG_H39<=zero;
XbG_H390<=zero;
XbG_H391<=zero;
XbG_H392<=zero;
XbG_H393<=zero;
XbG_H394<=zero;
XbG_H395<=zero;
XbG_H396<=zero;
XbG_H397<=zero;
XbG_H398<=zero;
XbG_H399<=zero;
XbG_H4<=zero;
XbG_H40<=zero;
XbG_H400<=zero;
XbG_H401<=zero;
XbG_H402<=zero;
XbG_H403<=zero;
XbG_H404<=zero;
XbG_H405<=zero;
XbG_H406<=zero;
XbG_H407<=zero;
XbG_H408<=zero;
XbG_H409<=zero;
XbG_H41<=zero;
XbG_H410<=zero;
XbG_H411<=zero;
XbG_H412<=zero;
XbG_H413<=zero;
XbG_H414<=zero;
XbG_H415<=zero;
XbG_H416<=zero;
XbG_H417<=zero;
XbG_H418<=zero;
XbG_H419<=zero;
XbG_H42<=zero;
XbG_H420<=zero;
XbG_H421<=zero;
XbG_H422<=zero;
XbG_H423<=zero;
XbG_H424<=zero;
XbG_H425<=zero;
XbG_H426<=zero;
XbG_H427<=zero;
XbG_H428<=zero;
XbG_H429<=zero;
XbG_H43<=zero;
XbG_H430<=zero;
XbG_H431<=zero;
XbG_H432<=zero;
XbG_H433<=zero;
XbG_H434<=zero;
XbG_H435<=zero;
XbG_H436<=zero;
XbG_H437<=zero;
XbG_H438<=zero;
XbG_H439<=zero;
XbG_H44<=zero;
XbG_H440<=zero;
XbG_H441<=zero;
XbG_H442<=zero;
XbG_H443<=zero;
XbG_H444<=zero;
XbG_H445<=zero;
XbG_H446<=zero;
XbG_H447<=zero;
XbG_H448<=zero;
XbG_H449<=zero;
XbG_H45<=zero;
XbG_H450<=zero;
XbG_H451<=zero;
XbG_H452<=zero;
XbG_H453<=zero;
XbG_H454<=zero;
XbG_H455<=zero;
XbG_H456<=zero;
XbG_H457<=zero;
XbG_H458<=zero;
XbG_H459<=zero;
XbG_H46<=zero;
XbG_H460<=zero;
XbG_H461<=zero;
XbG_H462<=zero;
XbG_H463<=zero;
XbG_H464<=zero;
XbG_H465<=zero;
XbG_H466<=zero;
XbG_H467<=zero;
XbG_H468<=zero;
XbG_H469<=zero;
XbG_H47<=zero;
XbG_H470<=zero;
XbG_H471<=zero;
XbG_H472<=zero;
XbG_H473<=zero;
XbG_H474<=zero;
XbG_H475<=zero;
XbG_H476<=zero;
XbG_H477<=zero;
XbG_H478<=zero;
XbG_H479<=zero;
XbG_H48<=zero;
XbG_H480<=zero;
XbG_H481<=zero;
XbG_H482<=zero;
XbG_H483<=zero;
XbG_H484<=zero;
XbG_H485<=zero;
XbG_H486<=zero;
XbG_H487<=zero;
XbG_H488<=zero;
XbG_H489<=zero;
XbG_H49<=zero;
XbG_H490<=zero;
XbG_H491<=zero;
XbG_H492<=zero;
XbG_H493<=zero;
XbG_H494<=zero;
XbG_H495<=zero;
XbG_H496<=zero;
XbG_H497<=zero;
XbG_H498<=zero;
XbG_H499<=zero;
XbG_H5<=zero;
XbG_H50<=zero;
XbG_H500<=zero;
XbG_H501<=zero;
XbG_H502<=zero;
XbG_H503<=zero;
XbG_H504<=zero;
XbG_H505<=zero;
XbG_H506<=zero;
XbG_H507<=zero;
XbG_H508<=zero;
XbG_H509<=zero;
XbG_H51<=zero;
XbG_H510<=zero;
XbG_H511<=zero;
XbG_H512<=zero;
XbG_H513<=zero;
XbG_H514<=zero;
XbG_H515<=zero;
XbG_H516<=zero;
XbG_H517<=zero;
XbG_H518<=zero;
XbG_H519<=zero;
XbG_H52<=zero;
XbG_H520<=zero;
XbG_H521<=zero;
XbG_H522<=zero;
XbG_H523<=zero;
XbG_H524<=zero;
XbG_H525<=zero;
XbG_H526<=zero;
XbG_H527<=zero;
XbG_H528<=zero;
XbG_H529<=zero;
XbG_H53<=zero;
XbG_H530<=zero;
XbG_H531<=zero;
XbG_H532<=zero;
XbG_H533<=zero;
XbG_H534<=zero;
XbG_H535<=zero;
XbG_H536<=zero;
XbG_H537<=zero;
XbG_H538<=zero;
XbG_H539<=zero;
XbG_H54<=zero;
XbG_H540<=zero;
XbG_H541<=zero;
XbG_H542<=zero;
XbG_H543<=zero;
XbG_H544<=zero;
XbG_H545<=zero;
XbG_H546<=zero;
XbG_H547<=zero;
XbG_H548<=zero;
XbG_H549<=zero;
XbG_H55<=zero;
XbG_H550<=zero;
XbG_H551<=zero;
XbG_H552<=zero;
XbG_H553<=zero;
XbG_H554<=zero;
XbG_H555<=zero;
XbG_H556<=zero;
XbG_H557<=zero;
XbG_H558<=zero;
XbG_H559<=zero;
XbG_H56<=zero;
XbG_H560<=zero;
XbG_H561<=zero;
XbG_H562<=zero;
XbG_H563<=zero;
XbG_H564<=zero;
XbG_H565<=zero;
XbG_H566<=zero;
XbG_H567<=zero;
XbG_H568<=zero;
XbG_H569<=zero;
XbG_H57<=zero;
XbG_H570<=zero;
XbG_H571<=zero;
XbG_H572<=zero;
XbG_H573<=zero;
XbG_H574<=zero;
XbG_H575<=zero;
XbG_H576<=zero;
XbG_H577<=zero;
XbG_H578<=zero;
XbG_H579<=zero;
XbG_H58<=zero;
XbG_H580<=zero;
XbG_H581<=zero;
XbG_H582<=zero;
XbG_H583<=zero;
XbG_H584<=zero;
XbG_H585<=zero;
XbG_H586<=zero;
XbG_H587<=zero;
XbG_H588<=zero;
XbG_H589<=zero;
XbG_H59<=zero;
XbG_H590<=zero;
XbG_H591<=zero;
XbG_H592<=zero;
XbG_H593<=zero;
XbG_H594<=zero;
XbG_H595<=zero;
XbG_H596<=zero;
XbG_H597<=zero;
XbG_H598<=zero;
XbG_H599<=zero;
XbG_H6<=zero;
XbG_H60<=zero;
XbG_H600<=zero;
XbG_H601<=zero;
XbG_H602<=zero;
XbG_H603<=zero;
XbG_H604<=zero;
XbG_H605<=zero;
XbG_H606<=zero;
XbG_H607<=zero;
XbG_H608<=zero;
XbG_H609<=zero;
XbG_H61<=zero;
XbG_H610<=zero;
XbG_H611<=zero;
XbG_H612<=zero;
XbG_H613<=zero;
XbG_H614<=zero;
XbG_H615<=zero;
XbG_H616<=zero;
XbG_H617<=zero;
XbG_H618<=zero;
XbG_H619<=zero;
XbG_H62<=zero;
XbG_H620<=zero;
XbG_H621<=zero;
XbG_H622<=zero;
XbG_H623<=zero;
XbG_H624<=zero;
XbG_H625<=zero;
XbG_H626<=zero;
XbG_H627<=zero;
XbG_H628<=zero;
XbG_H629<=zero;
XbG_H63<=zero;
XbG_H630<=zero;
XbG_H631<=zero;
XbG_H632<=zero;
XbG_H633<=zero;
XbG_H634<=zero;
XbG_H635<=zero;
XbG_H636<=zero;
XbG_H637<=zero;
XbG_H638<=zero;
XbG_H639<=zero;
XbG_H64<=zero;
XbG_H640<=zero;
XbG_H641<=zero;
XbG_H642<=zero;
XbG_H643<=zero;
XbG_H644<=zero;
XbG_H645<=zero;
XbG_H646<=zero;
XbG_H647<=zero;
XbG_H648<=zero;
XbG_H649<=zero;
XbG_H65<=zero;
XbG_H650<=zero;
XbG_H651<=zero;
XbG_H652<=zero;
XbG_H653<=zero;
XbG_H654<=zero;
XbG_H655<=zero;
XbG_H656<=zero;
XbG_H657<=zero;
XbG_H658<=zero;
XbG_H659<=zero;
XbG_H66<=zero;
XbG_H660<=zero;
XbG_H661<=Vr;
XbG_H662<=Vr;
XbG_H663<=Vr;
XbG_H664<=Vr;
XbG_H665<=Vr;
XbG_H666<=Vr;
XbG_H667<=Vr;
XbG_H668<=Vr;
XbG_H669<=Vr;
XbG_H67<=zero;
XbG_H670<=Vr;
XbG_H671<=Vr;
XbG_H672<=Vr;
XbG_H673<=Vr;
XbG_H674<=Vr;
XbG_H675<=Vr;
XbG_H676<=Vr;
XbG_H677<=Vr;
XbG_H678<=Vr;
XbG_H679<=Vr;
XbG_H68<=zero;
XbG_H680<=Vr;
XbG_H681<=Vr;
XbG_H682<=Vr;
XbG_H683<=Vr;
XbG_H684<=Vr;
XbG_H685<=Vr;
XbG_H686<=Vr;
XbG_H687<=Vr;
XbG_H688<=Vr;
XbG_H689<=Vr;
XbG_H69<=zero;
XbG_H690<=Vr;
XbG_H691<=Vr;
XbG_H692<=Vr;
XbG_H693<=Vr;
XbG_H694<=Vr;
XbG_H695<=Vr;
XbG_H696<=Vr;
XbG_H697<=Vr;
XbG_H698<=Vr;
XbG_H699<=Vr;
XbG_H7<=zero;
XbG_H70<=zero;
XbG_H700<=Vr;
XbG_H701<=Vr;
XbG_H702<=Vr;
XbG_H703<=Vr;
XbG_H704<=Vr;
XbG_H705<=Vr;
XbG_H706<=Vr;
XbG_H707<=Vr;
XbG_H708<=Vr;
XbG_H709<=Vr;
XbG_H71<=zero;
XbG_H710<=Vr;
XbG_H711<=Vr;
XbG_H712<=Vr;
XbG_H713<=Vr;
XbG_H714<=Vr;
XbG_H715<=Vr;
XbG_H716<=Vr;
XbG_H717<=Vr;
XbG_H718<=Vr;
XbG_H719<=Vr;
XbG_H72<=zero;
XbG_H720<=Vr;
XbG_H721<=Vr;
XbG_H722<=Vw;
XbG_H723<=Vw;
XbG_H724<=Vw;
XbG_H725<=Vw;
XbG_H726<=Vw;
XbG_H727<=Vw;
XbG_H728<=Vw;
XbG_H729<=Vw;
XbG_H73<=zero;
XbG_H730<=Vw;
XbG_H731<=Vw;
XbG_H732<=Vw;
XbG_H733<=Vw;
XbG_H734<=Vw;
XbG_H735<=Vw;
XbG_H74<=zero;
XbG_H75<=zero;
XbG_H76<=zero;
XbG_H77<=zero;
XbG_H78<=zero;
XbG_H79<=zero;
XbG_H8<=zero;
XbG_H80<=zero;
XbG_H81<=zero;
XbG_H82<=zero;
XbG_H83<=zero;
XbG_H84<=zero;
XbG_H85<=zero;
XbG_H86<=zero;
XbG_H87<=zero;
XbG_H88<=zero;
XbG_H89<=zero;
XbG_H9<=zero;
XbG_H90<=zero;
XbG_H91<=zero;
XbG_H92<=zero;
XbG_H93<=zero;
XbG_H94<=zero;
XbG_H95<=zero;
XbG_H96<=zero;
XbG_H97<=zero;
XbG_H98<=zero;
XbG_H99<=zero;
XbG_V0<=(others=>'Z');
XbG_V1<=(others=>'Z');
XbG_V10<=Vr, (others=>'Z') after 1 ps;
XbG_V100<=Vr;
XbG_V101<=Vr;
XbG_V102<=Vr;
XbG_V103<=Vr;
XbG_V104<=Vr;
XbG_V105<=Vr;
XbG_V106<=Vr;
XbG_V107<=Vr;
XbG_V108<=Vr;
XbG_V109<=Vr;
XbG_V11<=Vr, (others=>'Z') after 1 ps;
XbG_V110<=Vr;
XbG_V111<=Vr;
XbG_V112<=Vr;
XbG_V113<=Vr;
XbG_V114<=Vr;
XbG_V115<=Vr;
XbG_V116<=Vr;
XbG_V117<=Vr;
XbG_V118<=Vr;
XbG_V119<=Vr;
XbG_V12<=Vr, (others=>'Z') after 1 ps;
XbG_V120<=Vr;
XbG_V121<=Vr;
XbG_V122<=Vr;
XbG_V123<=Vr;
XbG_V124<=Vr;
XbG_V125<=Vr;
XbG_V126<=Vr;
XbG_V127<=Vr;
XbG_V128<=Vr;
XbG_V129<=Vr;
XbG_V13<=Vr, (others=>'Z') after 1 ps;
XbG_V130<=Vr;
XbG_V131<=Vr;
XbG_V132<=Vr;
XbG_V133<=Vr;
XbG_V134<=Vr;
XbG_V135<=Vr;
XbG_V136<=Vr;
XbG_V137<=Vr;
XbG_V138<=Vr;
XbG_V139<=Vr;
XbG_V14<=Vr, (others=>'Z') after 1 ps;
XbG_V140<=Vr;
XbG_V141<=Vr;
XbG_V142<=Vr;
XbG_V143<=Vr;
XbG_V144<=Vr;
XbG_V145<=Vr;
XbG_V146<=Vr;
XbG_V147<=Vr;
XbG_V148<=Vr;
XbG_V149<=Vr;
XbG_V15<=Vr, (others=>'Z') after 1 ps;
XbG_V150<=Vr;
XbG_V151<=Vr;
XbG_V152<=Vr;
XbG_V153<=Vr;
XbG_V154<=Vr;
XbG_V155<=Vr;
XbG_V156<=Vr;
XbG_V157<=Vr;
XbG_V158<=Vr;
XbG_V159<=Vr;
XbG_V16<=Vr, (others=>'Z') after 1 ps;
XbG_V160<=Vr;
XbG_V161<=Vr;
XbG_V162<=Vr;
XbG_V163<=Vr;
XbG_V164<=Vr;
XbG_V165<=Vr;
XbG_V166<=Vr;
XbG_V167<=Vr;
XbG_V168<=Vr;
XbG_V169<=Vr;
XbG_V17<=Vr, (others=>'Z') after 1 ps;
XbG_V170<=Vr;
XbG_V171<=Vr;
XbG_V172<=Vr;
XbG_V173<=Vr;
XbG_V174<=Vr;
XbG_V175<=Vr;
XbG_V176<=zero;
XbG_V177<=zero;
XbG_V178<=zero;
XbG_V179<=zero;
XbG_V18<=(others=>'Z');
XbG_V180<=zero;
XbG_V181<=zero;
XbG_V182<=zero;
XbG_V183<=zero;
XbG_V184<=zero;
XbG_V185<=zero;
XbG_V186<=zero;
XbG_V187<=zero;
XbG_V188<=zero;
XbG_V189<=zero;
XbG_V19<=(others=>'Z');
XbG_V2<=(others=>'Z');
XbG_V20<=(others=>'Z');
XbG_V21<=(others=>'Z');
XbG_V22<=(others=>'Z');
XbG_V23<=(others=>'Z');
XbG_V24<=(others=>'Z');
XbG_V25<=(others=>'Z');
XbG_V26<=(others=>'Z');
XbG_V27<=(others=>'Z');
XbG_V28<=(others=>'Z');
XbG_V29<=(others=>'Z');
XbG_V3<=(others=>'Z');
XbG_V30<=(others=>'Z');
XbG_V31<=(others=>'Z');
XbG_V32<=(others=>'Z');
XbG_V33<=(others=>'Z');
XbG_V34<=(others=>'Z');
XbG_V35<=(others=>'Z');
XbG_V36<=(others=>'Z');
XbG_V37<=(others=>'Z');
XbG_V38<=(others=>'Z');
XbG_V39<=(others=>'Z');
XbG_V4<=Vr, (others=>'Z') after 1 ps;
XbG_V40<=(others=>'Z');
XbG_V41<=(others=>'Z');
XbG_V42<=(others=>'Z');
XbG_V43<=(others=>'Z');
XbG_V44<=(others=>'Z');
XbG_V45<=(others=>'Z');
XbG_V46<=(others=>'Z');
XbG_V47<=(others=>'Z');
XbG_V48<=(others=>'Z');
XbG_V49<=(others=>'Z');
XbG_V5<=Vr, (others=>'Z') after 1 ps;
XbG_V50<=(others=>'Z');
XbG_V51<=(others=>'Z');
XbG_V52<=(others=>'Z');
XbG_V53<=(others=>'Z');
XbG_V54<=(others=>'Z');
XbG_V55<=(others=>'Z');
XbG_V56<=(others=>'Z');
XbG_V57<=(others=>'Z');
XbG_V58<=(others=>'Z');
XbG_V59<=(others=>'Z');
XbG_V6<=Vr, (others=>'Z') after 1 ps;
XbG_V60<=(others=>'Z');
XbG_V61<=(others=>'Z');
XbG_V62<=(others=>'Z');
XbG_V63<=(others=>'Z');
XbG_V64<=(others=>'Z');
XbG_V65<=(others=>'Z');
XbG_V66<=(others=>'Z');
XbG_V67<=(others=>'Z');
XbG_V68<=Vr;
XbG_V69<=Vr;
XbG_V7<=Vr, (others=>'Z') after 1 ps;
XbG_V70<=Vr;
XbG_V71<=Vr;
XbG_V72<=Vr;
XbG_V73<=Vr;
XbG_V74<=Vr;
XbG_V75<=Vr;
XbG_V76<=Vr;
XbG_V77<=Vr;
XbG_V78<=Vr;
XbG_V79<=Vr;
XbG_V8<=Vr, (others=>'Z') after 1 ps;
XbG_V80<=Vr;
XbG_V81<=Vr;
XbG_V82<=Vr;
XbG_V83<=Vr;
XbG_V84<=Vr;
XbG_V85<=Vr;
XbG_V86<=Vr;
XbG_V87<=Vr;
XbG_V88<=Vr;
XbG_V89<=Vr;
XbG_V9<=Vr, (others=>'Z') after 1 ps;
XbG_V90<=Vr;
XbG_V91<=Vr;
XbG_V92<=Vr;
XbG_V93<=Vr;
XbG_V94<=Vr;
XbG_V95<=Vr;
XbG_V96<=Vr;
XbG_V97<=Vr;
XbG_V98<=Vr;
XbG_V99<=Vr;

next_state<=D_EVM;

when D_EVM =>

XbG_H0<=Vr;
XbG_H1<=(others=>'Z');
XbG_H10<=(others=>'Z');
XbG_H100<=(others=>'Z');
XbG_H101<=(others=>'Z');
XbG_H102<=(others=>'Z');
XbG_H103<=(others=>'Z');
XbG_H104<=(others=>'Z');
XbG_H105<=(others=>'Z');
XbG_H106<=(others=>'Z');
XbG_H107<=(others=>'Z');
XbG_H108<=(others=>'Z');
XbG_H109<=(others=>'Z');
XbG_H11<=(others=>'Z');
XbG_H110<=(others=>'Z');
XbG_H111<=(others=>'Z');
XbG_H112<=(others=>'Z');
XbG_H113<=(others=>'Z');
XbG_H114<=(others=>'Z');
XbG_H115<=(others=>'Z');
XbG_H116<=(others=>'Z');
XbG_H117<=(others=>'Z');
XbG_H118<=(others=>'Z');
XbG_H119<=(others=>'Z');
XbG_H12<=(others=>'Z');
XbG_H120<=(others=>'Z');
XbG_H121<=(others=>'Z');
XbG_H122<=(others=>'Z');
XbG_H123<=(others=>'Z');
XbG_H124<=(others=>'Z');
XbG_H125<=(others=>'Z');
XbG_H126<=(others=>'Z');
XbG_H127<=(others=>'Z');
XbG_H128<=(others=>'Z');
XbG_H129<=(others=>'Z');
XbG_H13<=(others=>'Z');
XbG_H130<=(others=>'Z');
XbG_H131<=(others=>'Z');
XbG_H132<=(others=>'Z');
XbG_H133<=(others=>'Z');
XbG_H134<=(others=>'Z');
XbG_H135<=(others=>'Z');
XbG_H136<=(others=>'Z');
XbG_H137<=(others=>'Z');
XbG_H138<=(others=>'Z');
XbG_H139<=(others=>'Z');
XbG_H14<=(others=>'Z');
XbG_H140<=(others=>'Z');
XbG_H141<=(others=>'Z');
XbG_H142<=(others=>'Z');
XbG_H143<=(others=>'Z');
XbG_H144<=(others=>'Z');
XbG_H145<=(others=>'Z');
XbG_H146<=(others=>'Z');
XbG_H147<=(others=>'Z');
XbG_H148<=(others=>'Z');
XbG_H149<=(others=>'Z');
XbG_H15<=(others=>'Z');
XbG_H150<=(others=>'Z');
XbG_H151<=(others=>'Z');
XbG_H152<=(others=>'Z');
XbG_H153<=(others=>'Z');
XbG_H154<=(others=>'Z');
XbG_H155<=(others=>'Z');
XbG_H156<=(others=>'Z');
XbG_H157<=(others=>'Z');
XbG_H158<=(others=>'Z');
XbG_H159<=(others=>'Z');
XbG_H16<=(others=>'Z');
XbG_H160<=(others=>'Z');
XbG_H161<=(others=>'Z');
XbG_H162<=(others=>'Z');
XbG_H163<=(others=>'Z');
XbG_H164<=(others=>'Z');
XbG_H165<=(others=>'Z');
XbG_H166<=(others=>'Z');
XbG_H167<=(others=>'Z');
XbG_H168<=(others=>'Z');
XbG_H169<=(others=>'Z');
XbG_H17<=(others=>'Z');
XbG_H170<=(others=>'Z');
XbG_H171<=(others=>'Z');
XbG_H172<=(others=>'Z');
XbG_H173<=(others=>'Z');
XbG_H174<=(others=>'Z');
XbG_H175<=(others=>'Z');
XbG_H176<=(others=>'Z');
XbG_H177<=(others=>'Z');
XbG_H178<=(others=>'Z');
XbG_H179<=(others=>'Z');
XbG_H18<=(others=>'Z');
XbG_H180<=(others=>'Z');
XbG_H181<=(others=>'Z');
XbG_H182<=(others=>'Z');
XbG_H183<=(others=>'Z');
XbG_H184<=(others=>'Z');
XbG_H185<=(others=>'Z');
XbG_H186<=(others=>'Z');
XbG_H187<=(others=>'Z');
XbG_H188<=(others=>'Z');
XbG_H189<=(others=>'Z');
XbG_H19<=(others=>'Z');
XbG_H190<=(others=>'Z');
XbG_H191<=(others=>'Z');
XbG_H192<=(others=>'Z');
XbG_H193<=(others=>'Z');
XbG_H194<=(others=>'Z');
XbG_H195<=(others=>'Z');
XbG_H196<=(others=>'Z');
XbG_H197<=(others=>'Z');
XbG_H198<=(others=>'Z');
XbG_H199<=(others=>'Z');
XbG_H2<=(others=>'Z');
XbG_H20<=(others=>'Z');
XbG_H200<=(others=>'Z');
XbG_H201<=(others=>'Z');
XbG_H202<=(others=>'Z');
XbG_H203<=(others=>'Z');
XbG_H204<=(others=>'Z');
XbG_H205<=(others=>'Z');
XbG_H206<=(others=>'Z');
XbG_H207<=(others=>'Z');
XbG_H208<=(others=>'Z');
XbG_H209<=(others=>'Z');
XbG_H21<=(others=>'Z');
XbG_H210<=(others=>'Z');
XbG_H211<=(others=>'Z');
XbG_H212<=(others=>'Z');
XbG_H213<=(others=>'Z');
XbG_H214<=(others=>'Z');
XbG_H215<=(others=>'Z');
XbG_H216<=(others=>'Z');
XbG_H217<=(others=>'Z');
XbG_H218<=(others=>'Z');
XbG_H219<=(others=>'Z');
XbG_H22<=(others=>'Z');
XbG_H220<=(others=>'Z');
XbG_H221<=(others=>'Z');
XbG_H222<=(others=>'Z');
XbG_H223<=(others=>'Z');
XbG_H224<=(others=>'Z');
XbG_H225<=(others=>'Z');
XbG_H226<=(others=>'Z');
XbG_H227<=(others=>'Z');
XbG_H228<=(others=>'Z');
XbG_H229<=(others=>'Z');
XbG_H23<=(others=>'Z');
XbG_H230<=(others=>'Z');
XbG_H231<=(others=>'Z');
XbG_H232<=(others=>'Z');
XbG_H233<=(others=>'Z');
XbG_H234<=(others=>'Z');
XbG_H235<=(others=>'Z');
XbG_H236<=(others=>'Z');
XbG_H237<=(others=>'Z');
XbG_H238<=(others=>'Z');
XbG_H239<=(others=>'Z');
XbG_H24<=(others=>'Z');
XbG_H240<=(others=>'Z');
XbG_H241<=(others=>'Z');
XbG_H242<=(others=>'Z');
XbG_H243<=(others=>'Z');
XbG_H244<=(others=>'Z');
XbG_H245<=(others=>'Z');
XbG_H246<=(others=>'Z');
XbG_H247<=(others=>'Z');
XbG_H248<=(others=>'Z');
XbG_H249<=(others=>'Z');
XbG_H25<=(others=>'Z');
XbG_H250<=(others=>'Z');
XbG_H251<=(others=>'Z');
XbG_H252<=(others=>'Z');
XbG_H253<=(others=>'Z');
XbG_H254<=(others=>'Z');
XbG_H255<=(others=>'Z');
XbG_H256<=(others=>'Z');
XbG_H257<=(others=>'Z');
XbG_H258<=(others=>'Z');
XbG_H259<=(others=>'Z');
XbG_H26<=(others=>'Z');
XbG_H260<=(others=>'Z');
XbG_H261<=(others=>'Z');
XbG_H262<=(others=>'Z');
XbG_H263<=(others=>'Z');
XbG_H264<=(others=>'Z');
XbG_H265<=(others=>'Z');
XbG_H266<=(others=>'Z');
XbG_H267<=(others=>'Z');
XbG_H268<=(others=>'Z');
XbG_H269<=(others=>'Z');
XbG_H27<=(others=>'Z');
XbG_H270<=(others=>'Z');
XbG_H271<=(others=>'Z');
XbG_H272<=(others=>'Z');
XbG_H273<=(others=>'Z');
XbG_H274<=(others=>'Z');
XbG_H275<=(others=>'Z');
XbG_H276<=(others=>'Z');
XbG_H277<=(others=>'Z');
XbG_H278<=(others=>'Z');
XbG_H279<=(others=>'Z');
XbG_H28<=(others=>'Z');
XbG_H280<=(others=>'Z');
XbG_H281<=(others=>'Z');
XbG_H282<=(others=>'Z');
XbG_H283<=(others=>'Z');
XbG_H284<=(others=>'Z');
XbG_H285<=(others=>'Z');
XbG_H286<=(others=>'Z');
XbG_H287<=(others=>'Z');
XbG_H288<=(others=>'Z');
XbG_H289<=(others=>'Z');
XbG_H29<=(others=>'Z');
XbG_H290<=(others=>'Z');
XbG_H291<=(others=>'Z');
XbG_H292<=(others=>'Z');
XbG_H293<=(others=>'Z');
XbG_H294<=(others=>'Z');
XbG_H295<=(others=>'Z');
XbG_H296<=(others=>'Z');
XbG_H297<=(others=>'Z');
XbG_H298<=(others=>'Z');
XbG_H299<=(others=>'Z');
XbG_H3<=(others=>'Z');
XbG_H30<=(others=>'Z');
XbG_H300<=(others=>'Z');
XbG_H301<=(others=>'Z');
XbG_H302<=(others=>'Z');
XbG_H303<=(others=>'Z');
XbG_H304<=(others=>'Z');
XbG_H305<=(others=>'Z');
XbG_H306<=(others=>'Z');
XbG_H307<=(others=>'Z');
XbG_H308<=(others=>'Z');
XbG_H309<=(others=>'Z');
XbG_H31<=(others=>'Z');
XbG_H310<=(others=>'Z');
XbG_H311<=(others=>'Z');
XbG_H312<=(others=>'Z');
XbG_H313<=(others=>'Z');
XbG_H314<=(others=>'Z');
XbG_H315<=(others=>'Z');
XbG_H316<=(others=>'Z');
XbG_H317<=(others=>'Z');
XbG_H318<=(others=>'Z');
XbG_H319<=(others=>'Z');
XbG_H32<=(others=>'Z');
XbG_H320<=(others=>'Z');
XbG_H321<=(others=>'Z');
XbG_H322<=(others=>'Z');
XbG_H323<=(others=>'Z');
XbG_H324<=(others=>'Z');
XbG_H325<=(others=>'Z');
XbG_H326<=(others=>'Z');
XbG_H327<=(others=>'Z');
XbG_H328<=(others=>'Z');
XbG_H329<=(others=>'Z');
XbG_H33<=(others=>'Z');
XbG_H330<=(others=>'Z');
XbG_H331<=(others=>'Z');
XbG_H332<=(others=>'Z');
XbG_H333<=(others=>'Z');
XbG_H334<=(others=>'Z');
XbG_H335<=(others=>'Z');
XbG_H336<=(others=>'Z');
XbG_H337<=(others=>'Z');
XbG_H338<=(others=>'Z');
XbG_H339<=(others=>'Z');
XbG_H34<=(others=>'Z');
XbG_H340<=(others=>'Z');
XbG_H341<=(others=>'Z');
XbG_H342<=(others=>'Z');
XbG_H343<=(others=>'Z');
XbG_H344<=(others=>'Z');
XbG_H345<=(others=>'Z');
XbG_H346<=(others=>'Z');
XbG_H347<=(others=>'Z');
XbG_H348<=(others=>'Z');
XbG_H349<=(others=>'Z');
XbG_H35<=(others=>'Z');
XbG_H350<=(others=>'Z');
XbG_H351<=(others=>'Z');
XbG_H352<=(others=>'Z');
XbG_H353<=(others=>'Z');
XbG_H354<=(others=>'Z');
XbG_H355<=(others=>'Z');
XbG_H356<=(others=>'Z');
XbG_H357<=(others=>'Z');
XbG_H358<=(others=>'Z');
XbG_H359<=(others=>'Z');
XbG_H36<=(others=>'Z');
XbG_H360<=(others=>'Z');
XbG_H361<=(others=>'Z');
XbG_H362<=(others=>'Z');
XbG_H363<=(others=>'Z');
XbG_H364<=(others=>'Z');
XbG_H365<=(others=>'Z');
XbG_H366<=(others=>'Z');
XbG_H367<=(others=>'Z');
XbG_H368<=(others=>'Z');
XbG_H369<=(others=>'Z');
XbG_H37<=(others=>'Z');
XbG_H370<=(others=>'Z');
XbG_H371<=(others=>'Z');
XbG_H372<=(others=>'Z');
XbG_H373<=(others=>'Z');
XbG_H374<=(others=>'Z');
XbG_H375<=(others=>'Z');
XbG_H376<=(others=>'Z');
XbG_H377<=(others=>'Z');
XbG_H378<=(others=>'Z');
XbG_H379<=(others=>'Z');
XbG_H38<=(others=>'Z');
XbG_H380<=(others=>'Z');
XbG_H381<=(others=>'Z');
XbG_H382<=(others=>'Z');
XbG_H383<=(others=>'Z');
XbG_H384<=(others=>'Z');
XbG_H385<=(others=>'Z');
XbG_H386<=(others=>'Z');
XbG_H387<=(others=>'Z');
XbG_H388<=(others=>'Z');
XbG_H389<=(others=>'Z');
XbG_H39<=(others=>'Z');
XbG_H390<=(others=>'Z');
XbG_H391<=(others=>'Z');
XbG_H392<=(others=>'Z');
XbG_H393<=(others=>'Z');
XbG_H394<=(others=>'Z');
XbG_H395<=(others=>'Z');
XbG_H396<=(others=>'Z');
XbG_H397<=(others=>'Z');
XbG_H398<=(others=>'Z');
XbG_H399<=(others=>'Z');
XbG_H4<=(others=>'Z');
XbG_H40<=(others=>'Z');
XbG_H400<=(others=>'Z');
XbG_H401<=(others=>'Z');
XbG_H402<=(others=>'Z');
XbG_H403<=(others=>'Z');
XbG_H404<=(others=>'Z');
XbG_H405<=(others=>'Z');
XbG_H406<=(others=>'Z');
XbG_H407<=(others=>'Z');
XbG_H408<=(others=>'Z');
XbG_H409<=(others=>'Z');
XbG_H41<=(others=>'Z');
XbG_H410<=(others=>'Z');
XbG_H411<=(others=>'Z');
XbG_H412<=(others=>'Z');
XbG_H413<=(others=>'Z');
XbG_H414<=(others=>'Z');
XbG_H415<=(others=>'Z');
XbG_H416<=(others=>'Z');
XbG_H417<=(others=>'Z');
XbG_H418<=(others=>'Z');
XbG_H419<=(others=>'Z');
XbG_H42<=(others=>'Z');
XbG_H420<=(others=>'Z');
XbG_H421<=(others=>'Z');
XbG_H422<=(others=>'Z');
XbG_H423<=(others=>'Z');
XbG_H424<=(others=>'Z');
XbG_H425<=(others=>'Z');
XbG_H426<=(others=>'Z');
XbG_H427<=(others=>'Z');
XbG_H428<=(others=>'Z');
XbG_H429<=(others=>'Z');
XbG_H43<=(others=>'Z');
XbG_H430<=(others=>'Z');
XbG_H431<=(others=>'Z');
XbG_H432<=(others=>'Z');
XbG_H433<=(others=>'Z');
XbG_H434<=(others=>'Z');
XbG_H435<=(others=>'Z');
XbG_H436<=(others=>'Z');
XbG_H437<=(others=>'Z');
XbG_H438<=(others=>'Z');
XbG_H439<=(others=>'Z');
XbG_H44<=(others=>'Z');
XbG_H440<=(others=>'Z');
XbG_H441<=(others=>'Z');
XbG_H442<=(others=>'Z');
XbG_H443<=(others=>'Z');
XbG_H444<=(others=>'Z');
XbG_H445<=(others=>'Z');
XbG_H446<=(others=>'Z');
XbG_H447<=(others=>'Z');
XbG_H448<=(others=>'Z');
XbG_H449<=(others=>'Z');
XbG_H45<=(others=>'Z');
XbG_H450<=(others=>'Z');
XbG_H451<=(others=>'Z');
XbG_H452<=(others=>'Z');
XbG_H453<=(others=>'Z');
XbG_H454<=(others=>'Z');
XbG_H455<=(others=>'Z');
XbG_H456<=(others=>'Z');
XbG_H457<=(others=>'Z');
XbG_H458<=(others=>'Z');
XbG_H459<=(others=>'Z');
XbG_H46<=(others=>'Z');
XbG_H460<=(others=>'Z');
XbG_H461<=(others=>'Z');
XbG_H462<=(others=>'Z');
XbG_H463<=(others=>'Z');
XbG_H464<=(others=>'Z');
XbG_H465<=(others=>'Z');
XbG_H466<=(others=>'Z');
XbG_H467<=(others=>'Z');
XbG_H468<=(others=>'Z');
XbG_H469<=(others=>'Z');
XbG_H47<=(others=>'Z');
XbG_H470<=(others=>'Z');
XbG_H471<=(others=>'Z');
XbG_H472<=(others=>'Z');
XbG_H473<=(others=>'Z');
XbG_H474<=(others=>'Z');
XbG_H475<=(others=>'Z');
XbG_H476<=(others=>'Z');
XbG_H477<=(others=>'Z');
XbG_H478<=(others=>'Z');
XbG_H479<=(others=>'Z');
XbG_H48<=(others=>'Z');
XbG_H480<=(others=>'Z');
XbG_H481<=(others=>'Z');
XbG_H482<=(others=>'Z');
XbG_H483<=(others=>'Z');
XbG_H484<=(others=>'Z');
XbG_H485<=(others=>'Z');
XbG_H486<=(others=>'Z');
XbG_H487<=(others=>'Z');
XbG_H488<=(others=>'Z');
XbG_H489<=(others=>'Z');
XbG_H49<=(others=>'Z');
XbG_H490<=(others=>'Z');
XbG_H491<=(others=>'Z');
XbG_H492<=(others=>'Z');
XbG_H493<=(others=>'Z');
XbG_H494<=(others=>'Z');
XbG_H495<=(others=>'Z');
XbG_H496<=(others=>'Z');
XbG_H497<=(others=>'Z');
XbG_H498<=(others=>'Z');
XbG_H499<=(others=>'Z');
XbG_H5<=(others=>'Z');
XbG_H50<=(others=>'Z');
XbG_H500<=(others=>'Z');
XbG_H501<=(others=>'Z');
XbG_H502<=(others=>'Z');
XbG_H503<=(others=>'Z');
XbG_H504<=(others=>'Z');
XbG_H505<=(others=>'Z');
XbG_H506<=(others=>'Z');
XbG_H507<=(others=>'Z');
XbG_H508<=(others=>'Z');
XbG_H509<=(others=>'Z');
XbG_H51<=(others=>'Z');
XbG_H510<=(others=>'Z');
XbG_H511<=(others=>'Z');
XbG_H512<=(others=>'Z');
XbG_H513<=(others=>'Z');
XbG_H514<=(others=>'Z');
XbG_H515<=(others=>'Z');
XbG_H516<=(others=>'Z');
XbG_H517<=(others=>'Z');
XbG_H518<=(others=>'Z');
XbG_H519<=(others=>'Z');
XbG_H52<=(others=>'Z');
XbG_H520<=(others=>'Z');
XbG_H521<=(others=>'Z');
XbG_H522<=(others=>'Z');
XbG_H523<=(others=>'Z');
XbG_H524<=(others=>'Z');
XbG_H525<=(others=>'Z');
XbG_H526<=(others=>'Z');
XbG_H527<=(others=>'Z');
XbG_H528<=(others=>'Z');
XbG_H529<=(others=>'Z');
XbG_H53<=(others=>'Z');
XbG_H530<=(others=>'Z');
XbG_H531<=(others=>'Z');
XbG_H532<=(others=>'Z');
XbG_H533<=(others=>'Z');
XbG_H534<=(others=>'Z');
XbG_H535<=(others=>'Z');
XbG_H536<=(others=>'Z');
XbG_H537<=(others=>'Z');
XbG_H538<=(others=>'Z');
XbG_H539<=(others=>'Z');
XbG_H54<=(others=>'Z');
XbG_H540<=(others=>'Z');
XbG_H541<=(others=>'Z');
XbG_H542<=(others=>'Z');
XbG_H543<=(others=>'Z');
XbG_H544<=(others=>'Z');
XbG_H545<=(others=>'Z');
XbG_H546<=(others=>'Z');
XbG_H547<=(others=>'Z');
XbG_H548<=(others=>'Z');
XbG_H549<=(others=>'Z');
XbG_H55<=(others=>'Z');
XbG_H550<=(others=>'Z');
XbG_H551<=(others=>'Z');
XbG_H552<=(others=>'Z');
XbG_H553<=(others=>'Z');
XbG_H554<=(others=>'Z');
XbG_H555<=(others=>'Z');
XbG_H556<=(others=>'Z');
XbG_H557<=(others=>'Z');
XbG_H558<=(others=>'Z');
XbG_H559<=(others=>'Z');
XbG_H56<=(others=>'Z');
XbG_H560<=(others=>'Z');
XbG_H561<=(others=>'Z');
XbG_H562<=(others=>'Z');
XbG_H563<=(others=>'Z');
XbG_H564<=(others=>'Z');
XbG_H565<=(others=>'Z');
XbG_H566<=(others=>'Z');
XbG_H567<=(others=>'Z');
XbG_H568<=(others=>'Z');
XbG_H569<=(others=>'Z');
XbG_H57<=(others=>'Z');
XbG_H570<=(others=>'Z');
XbG_H571<=(others=>'Z');
XbG_H572<=(others=>'Z');
XbG_H573<=(others=>'Z');
XbG_H574<=(others=>'Z');
XbG_H575<=(others=>'Z');
XbG_H576<=(others=>'Z');
XbG_H577<=(others=>'Z');
XbG_H578<=(others=>'Z');
XbG_H579<=(others=>'Z');
XbG_H58<=(others=>'Z');
XbG_H580<=(others=>'Z');
XbG_H581<=(others=>'Z');
XbG_H582<=(others=>'Z');
XbG_H583<=(others=>'Z');
XbG_H584<=(others=>'Z');
XbG_H585<=(others=>'Z');
XbG_H586<=(others=>'Z');
XbG_H587<=(others=>'Z');
XbG_H588<=(others=>'Z');
XbG_H589<=(others=>'Z');
XbG_H59<=(others=>'Z');
XbG_H590<=(others=>'Z');
XbG_H591<=(others=>'Z');
XbG_H592<=(others=>'Z');
XbG_H593<=(others=>'Z');
XbG_H594<=(others=>'Z');
XbG_H595<=(others=>'Z');
XbG_H596<=(others=>'Z');
XbG_H597<=(others=>'Z');
XbG_H598<=(others=>'Z');
XbG_H599<=(others=>'Z');
XbG_H6<=(others=>'Z');
XbG_H60<=(others=>'Z');
XbG_H600<=(others=>'Z');
XbG_H601<=(others=>'Z');
XbG_H602<=(others=>'Z');
XbG_H603<=(others=>'Z');
XbG_H604<=(others=>'Z');
XbG_H605<=(others=>'Z');
XbG_H606<=(others=>'Z');
XbG_H607<=(others=>'Z');
XbG_H608<=(others=>'Z');
XbG_H609<=(others=>'Z');
XbG_H61<=(others=>'Z');
XbG_H610<=(others=>'Z');
XbG_H611<=(others=>'Z');
XbG_H612<=(others=>'Z');
XbG_H613<=(others=>'Z');
XbG_H614<=(others=>'Z');
XbG_H615<=(others=>'Z');
XbG_H616<=(others=>'Z');
XbG_H617<=(others=>'Z');
XbG_H618<=(others=>'Z');
XbG_H619<=(others=>'Z');
XbG_H62<=(others=>'Z');
XbG_H620<=(others=>'Z');
XbG_H621<=(others=>'Z');
XbG_H622<=(others=>'Z');
XbG_H623<=(others=>'Z');
XbG_H624<=(others=>'Z');
XbG_H625<=(others=>'Z');
XbG_H626<=(others=>'Z');
XbG_H627<=(others=>'Z');
XbG_H628<=(others=>'Z');
XbG_H629<=(others=>'Z');
XbG_H63<=(others=>'Z');
XbG_H630<=(others=>'Z');
XbG_H631<=(others=>'Z');
XbG_H632<=(others=>'Z');
XbG_H633<=(others=>'Z');
XbG_H634<=(others=>'Z');
XbG_H635<=(others=>'Z');
XbG_H636<=(others=>'Z');
XbG_H637<=(others=>'Z');
XbG_H638<=(others=>'Z');
XbG_H639<=(others=>'Z');
XbG_H64<=(others=>'Z');
XbG_H640<=(others=>'Z');
XbG_H641<=(others=>'Z');
XbG_H642<=(others=>'Z');
XbG_H643<=(others=>'Z');
XbG_H644<=(others=>'Z');
XbG_H645<=(others=>'Z');
XbG_H646<=(others=>'Z');
XbG_H647<=(others=>'Z');
XbG_H648<=(others=>'Z');
XbG_H649<=(others=>'Z');
XbG_H65<=(others=>'Z');
XbG_H650<=(others=>'Z');
XbG_H651<=(others=>'Z');
XbG_H652<=(others=>'Z');
XbG_H653<=(others=>'Z');
XbG_H654<=(others=>'Z');
XbG_H655<=(others=>'Z');
XbG_H656<=(others=>'Z');
XbG_H657<=(others=>'Z');
XbG_H658<=(others=>'Z');
XbG_H659<=(others=>'Z');
XbG_H66<=(others=>'Z');
XbG_H660<=(others=>'Z');
XbG_H661<=Vr;
XbG_H662<=Vr;
XbG_H663<=Vr;
XbG_H664<=Vr;
XbG_H665<=Vr;
XbG_H666<=Vr;
XbG_H667<=Vr;
XbG_H668<=Vr;
XbG_H669<=Vr;
XbG_H67<=(others=>'Z');
XbG_H670<=Vr;
XbG_H671<=Vr;
XbG_H672<=Vr;
XbG_H673<=Vr;
XbG_H674<=Vr;
XbG_H675<=Vr;
XbG_H676<=Vr;
XbG_H677<=Vr;
XbG_H678<=Vr;
XbG_H679<=Vr;
XbG_H68<=(others=>'Z');
XbG_H680<=Vr;
XbG_H681<=Vr;
XbG_H682<=Vr;
XbG_H683<=Vr;
XbG_H684<=Vr;
XbG_H685<=Vr;
XbG_H686<=Vr;
XbG_H687<=Vr;
XbG_H688<=Vr;
XbG_H689<=Vr;
XbG_H69<=(others=>'Z');
XbG_H690<=Vr;
XbG_H691<=Vr;
XbG_H692<=Vr;
XbG_H693<=Vr;
XbG_H694<=Vr;
XbG_H695<=Vr;
XbG_H696<=Vr;
XbG_H697<=Vr;
XbG_H698<=Vr;
XbG_H699<=Vr;
XbG_H7<=(others=>'Z');
XbG_H70<=(others=>'Z');
XbG_H700<=Vr;
XbG_H701<=Vr;
XbG_H702<=Vr;
XbG_H703<=Vr;
XbG_H704<=Vr;
XbG_H705<=Vr;
XbG_H706<=Vr;
XbG_H707<=Vr;
XbG_H708<=Vr;
XbG_H709<=Vr;
XbG_H71<=(others=>'Z');
XbG_H710<=Vr;
XbG_H711<=Vr;
XbG_H712<=Vr;
XbG_H713<=Vr;
XbG_H714<=Vr;
XbG_H715<=Vr;
XbG_H716<=Vr;
XbG_H717<=Vr;
XbG_H718<=Vr;
XbG_H719<=Vr;
XbG_H72<=(others=>'Z');
XbG_H720<=Vr;
XbG_H721<=Vr;
XbG_H722<=Vr;
XbG_H723<=Vr;
XbG_H724<=Vr;
XbG_H725<=Vr;
XbG_H726<=Vr;
XbG_H727<=Vr;
XbG_H728<=Vr;
XbG_H729<=Vr;
XbG_H73<=(others=>'Z');
XbG_H730<=Vr;
XbG_H731<=Vr;
XbG_H732<=Vr;
XbG_H733<=Vr;
XbG_H734<=Vr;
XbG_H735<=Vr;
XbG_H74<=(others=>'Z');
XbG_H75<=(others=>'Z');
XbG_H76<=(others=>'Z');
XbG_H77<=(others=>'Z');
XbG_H78<=(others=>'Z');
XbG_H79<=(others=>'Z');
XbG_H8<=(others=>'Z');
XbG_H80<=(others=>'Z');
XbG_H81<=(others=>'Z');
XbG_H82<=(others=>'Z');
XbG_H83<=(others=>'Z');
XbG_H84<=(others=>'Z');
XbG_H85<=(others=>'Z');
XbG_H86<=(others=>'Z');
XbG_H87<=(others=>'Z');
XbG_H88<=(others=>'Z');
XbG_H89<=(others=>'Z');
XbG_H9<=(others=>'Z');
XbG_H90<=(others=>'Z');
XbG_H91<=(others=>'Z');
XbG_H92<=(others=>'Z');
XbG_H93<=(others=>'Z');
XbG_H94<=(others=>'Z');
XbG_H95<=(others=>'Z');
XbG_H96<=(others=>'Z');
XbG_H97<=(others=>'Z');
XbG_H98<=(others=>'Z');
XbG_H99<=(others=>'Z');
XbG_V0<=Vr;
XbG_V1<=Vr;
XbG_V10<=Vr;
XbG_V100<=Vr;
XbG_V101<=Vw;
XbG_V102<=Vr;
XbG_V103<=Vw;
XbG_V104<=Vr;
XbG_V105<=Vw;
XbG_V106<=Vr;
XbG_V107<=Vw;
XbG_V108<=Vr;
XbG_V109<=Vw;
XbG_V11<=Vr;
XbG_V110<=Vr;
XbG_V111<=Vw;
XbG_V112<=Vr;
XbG_V113<=Vw;
XbG_V114<=Vr;
XbG_V115<=Vw;
XbG_V116<=Vr;
XbG_V117<=Vw;
XbG_V118<=Vr;
XbG_V119<=Vw;
XbG_V12<=Vr;
XbG_V120<=Vr;
XbG_V121<=Vw;
XbG_V122<=Vr;
XbG_V123<=Vw;
XbG_V124<=Vr;
XbG_V125<=Vw;
XbG_V126<=Vr;
XbG_V127<=Vw;
XbG_V128<=Vr;
XbG_V129<=Vw;
XbG_V13<=Vr;
XbG_V130<=Vr;
XbG_V131<=Vw;
XbG_V132<=Vr;
XbG_V133<=Vw;
XbG_V134<=Vr;
XbG_V135<=Vw;
XbG_V136<=Vr;
XbG_V137<=Vw;
XbG_V138<=Vr;
XbG_V139<=Vw;
XbG_V14<=Vr;
XbG_V140<=Vr;
XbG_V141<=Vw;
XbG_V142<=Vr;
XbG_V143<=Vw;
XbG_V144<=Vr;
XbG_V145<=Vw;
XbG_V146<=Vr;
XbG_V147<=Vw;
XbG_V148<=Vr;
XbG_V149<=Vw;
XbG_V15<=Vr;
XbG_V150<=Vr;
XbG_V151<=Vw;
XbG_V152<=Vr;
XbG_V153<=Vw;
XbG_V154<=Vr;
XbG_V155<=Vw;
XbG_V156<=Vr;
XbG_V157<=Vw;
XbG_V158<=Vr;
XbG_V159<=Vw;
XbG_V16<=Vr;
XbG_V160<=Vr;
XbG_V161<=Vw;
XbG_V162<=Vr;
XbG_V163<=Vw;
XbG_V164<=Vr;
XbG_V165<=Vw;
XbG_V166<=Vr;
XbG_V167<=Vw;
XbG_V168<=Vr;
XbG_V169<=Vw;
XbG_V17<=Vr;
XbG_V170<=Vr;
XbG_V171<=Vw;
XbG_V172<=Vr;
XbG_V173<=Vw;
XbG_V174<=Vr;
XbG_V175<=Vw;
XbG_V176<=Vr;
XbG_V177<=Vw;
XbG_V178<=Vr;
XbG_V179<=Vw;
XbG_V18<=Vr;
XbG_V180<=Vr;
XbG_V181<=Vw;
XbG_V182<=Vr;
XbG_V183<=Vw;
XbG_V184<=Vr;
XbG_V185<=Vw;
XbG_V186<=Vr;
XbG_V187<=Vw;
XbG_V188<=Vr;
XbG_V189<=Vw;
XbG_V19<=Vr;
XbG_V2<=Vr;
XbG_V20<=Vr;
XbG_V21<=Vr;
XbG_V22<=Vr;
XbG_V23<=Vr;
XbG_V24<=Vr;
XbG_V25<=Vr;
XbG_V26<=Vr;
XbG_V27<=Vr;
XbG_V28<=Vr;
XbG_V29<=Vr;
XbG_V3<=Vr;
XbG_V30<=Vr;
XbG_V31<=Vr;
XbG_V32<=Vr;
XbG_V33<=Vr;
XbG_V34<=Vr;
XbG_V35<=Vr;
XbG_V36<=Vr;
XbG_V37<=Vr;
XbG_V38<=Vr;
XbG_V39<=Vr;
XbG_V4<=Vr;
XbG_V40<=Vr;
XbG_V41<=Vr;
XbG_V42<=Vr;
XbG_V43<=Vr;
XbG_V44<=Vr;
XbG_V45<=Vr;
XbG_V46<=Vr;
XbG_V47<=Vr;
XbG_V48<=Vr;
XbG_V49<=Vr;
XbG_V5<=Vr;
XbG_V50<=Vr;
XbG_V51<=Vr;
XbG_V52<=Vr;
XbG_V53<=Vr;
XbG_V54<=Vr;
XbG_V55<=Vr;
XbG_V56<=Vr;
XbG_V57<=Vr;
XbG_V58<=Vr;
XbG_V59<=Vr;
XbG_V6<=Vr;
XbG_V60<=Vr;
XbG_V61<=Vr;
XbG_V62<=Vr;
XbG_V63<=Vr;
XbG_V64<=Vr;
XbG_V65<=Vr;
XbG_V66<=Vr;
XbG_V67<=Vr;
XbG_V68<=Vr;
XbG_V69<=Vw;
XbG_V7<=Vr;
XbG_V70<=Vr;
XbG_V71<=Vw;
XbG_V72<=Vr;
XbG_V73<=Vw;
XbG_V74<=Vr;
XbG_V75<=Vw;
XbG_V76<=Vr;
XbG_V77<=Vw;
XbG_V78<=Vr;
XbG_V79<=Vw;
XbG_V8<=Vr;
XbG_V80<=Vr;
XbG_V81<=Vw;
XbG_V82<=Vr;
XbG_V83<=Vw;
XbG_V84<=Vr;
XbG_V85<=Vw;
XbG_V86<=Vr;
XbG_V87<=Vw;
XbG_V88<=Vr;
XbG_V89<=Vw;
XbG_V9<=Vr;
XbG_V90<=Vr;
XbG_V91<=Vw;
XbG_V92<=Vr;
XbG_V93<=Vw;
XbG_V94<=Vr;
XbG_V95<=Vw;
XbG_V96<=Vr;
XbG_V97<=Vw;
XbG_V98<=Vr;
XbG_V99<=Vw;

next_state<=E_EVR;

when E_EVR =>

XbG_H0<=Vr;
XbG_H1<=Vw;
XbG_H10<=Vw;
XbG_H100<=Vw;
XbG_H101<=Vw;
XbG_H102<=Vw;
XbG_H103<=Vw;
XbG_H104<=Vw;
XbG_H105<=Vw;
XbG_H106<=Vw;
XbG_H107<=Vw;
XbG_H108<=Vw;
XbG_H109<=Vw;
XbG_H11<=Vw;
XbG_H110<=Vw;
XbG_H111<=Vw;
XbG_H112<=Vw;
XbG_H113<=Vw;
XbG_H114<=Vw;
XbG_H115<=Vw;
XbG_H116<=Vw;
XbG_H117<=Vw;
XbG_H118<=Vw;
XbG_H119<=Vw;
XbG_H12<=Vw;
XbG_H120<=Vw;
XbG_H121<=Vw;
XbG_H122<=Vw;
XbG_H123<=Vw;
XbG_H124<=Vw;
XbG_H125<=Vw;
XbG_H126<=Vw;
XbG_H127<=Vw;
XbG_H128<=Vw;
XbG_H129<=Vw;
XbG_H13<=Vw;
XbG_H130<=Vw;
XbG_H131<=Vw;
XbG_H132<=Vw;
XbG_H133<=Vw;
XbG_H134<=Vw;
XbG_H135<=Vw;
XbG_H136<=Vw;
XbG_H137<=Vw;
XbG_H138<=Vw;
XbG_H139<=Vw;
XbG_H14<=Vw;
XbG_H140<=Vw;
XbG_H141<=Vw;
XbG_H142<=Vw;
XbG_H143<=Vw;
XbG_H144<=Vw;
XbG_H145<=Vw;
XbG_H146<=Vw;
XbG_H147<=Vw;
XbG_H148<=Vw;
XbG_H149<=Vw;
XbG_H15<=Vw;
XbG_H150<=Vw;
XbG_H151<=Vw;
XbG_H152<=Vw;
XbG_H153<=Vw;
XbG_H154<=Vw;
XbG_H155<=Vw;
XbG_H156<=Vw;
XbG_H157<=Vw;
XbG_H158<=Vw;
XbG_H159<=Vw;
XbG_H16<=Vw;
XbG_H160<=Vw;
XbG_H161<=Vw;
XbG_H162<=Vw;
XbG_H163<=Vw;
XbG_H164<=Vw;
XbG_H165<=Vw;
XbG_H166<=Vw;
XbG_H167<=Vw;
XbG_H168<=Vw;
XbG_H169<=Vw;
XbG_H17<=Vw;
XbG_H170<=Vw;
XbG_H171<=Vw;
XbG_H172<=Vw;
XbG_H173<=Vw;
XbG_H174<=Vw;
XbG_H175<=Vw;
XbG_H176<=Vw;
XbG_H177<=Vw;
XbG_H178<=Vw;
XbG_H179<=Vw;
XbG_H18<=Vw;
XbG_H180<=Vw;
XbG_H181<=Vw;
XbG_H182<=Vw;
XbG_H183<=Vw;
XbG_H184<=Vw;
XbG_H185<=Vw;
XbG_H186<=Vw;
XbG_H187<=Vw;
XbG_H188<=Vw;
XbG_H189<=Vw;
XbG_H19<=Vw;
XbG_H190<=Vw;
XbG_H191<=Vw;
XbG_H192<=Vw;
XbG_H193<=Vw;
XbG_H194<=Vw;
XbG_H195<=Vw;
XbG_H196<=Vw;
XbG_H197<=Vw;
XbG_H198<=Vw;
XbG_H199<=Vw;
XbG_H2<=Vw;
XbG_H20<=Vw;
XbG_H200<=Vw;
XbG_H201<=Vw;
XbG_H202<=Vw;
XbG_H203<=Vw;
XbG_H204<=Vw;
XbG_H205<=Vw;
XbG_H206<=Vw;
XbG_H207<=Vw;
XbG_H208<=Vw;
XbG_H209<=Vw;
XbG_H21<=Vw;
XbG_H210<=Vw;
XbG_H211<=Vw;
XbG_H212<=Vw;
XbG_H213<=Vw;
XbG_H214<=Vw;
XbG_H215<=Vw;
XbG_H216<=Vw;
XbG_H217<=Vw;
XbG_H218<=Vw;
XbG_H219<=Vw;
XbG_H22<=Vw;
XbG_H220<=Vw;
XbG_H221<=Vw;
XbG_H222<=Vw;
XbG_H223<=Vw;
XbG_H224<=Vw;
XbG_H225<=Vw;
XbG_H226<=Vw;
XbG_H227<=Vw;
XbG_H228<=Vw;
XbG_H229<=Vw;
XbG_H23<=Vw;
XbG_H230<=Vw;
XbG_H231<=Vw;
XbG_H232<=Vw;
XbG_H233<=Vw;
XbG_H234<=Vw;
XbG_H235<=Vw;
XbG_H236<=Vw;
XbG_H237<=Vw;
XbG_H238<=Vw;
XbG_H239<=Vw;
XbG_H24<=Vw;
XbG_H240<=Vw;
XbG_H241<=Vw;
XbG_H242<=Vw;
XbG_H243<=Vw;
XbG_H244<=Vw;
XbG_H245<=Vw;
XbG_H246<=Vw;
XbG_H247<=Vw;
XbG_H248<=Vw;
XbG_H249<=Vw;
XbG_H25<=Vw;
XbG_H250<=Vw;
XbG_H251<=Vw;
XbG_H252<=Vw;
XbG_H253<=Vw;
XbG_H254<=Vw;
XbG_H255<=Vw;
XbG_H256<=Vw;
XbG_H257<=Vw;
XbG_H258<=Vw;
XbG_H259<=Vw;
XbG_H26<=Vw;
XbG_H260<=Vw;
XbG_H261<=Vw;
XbG_H262<=Vw;
XbG_H263<=Vw;
XbG_H264<=Vw;
XbG_H265<=Vw;
XbG_H266<=Vw;
XbG_H267<=Vw;
XbG_H268<=Vw;
XbG_H269<=Vw;
XbG_H27<=Vw;
XbG_H270<=Vw;
XbG_H271<=Vw;
XbG_H272<=Vw;
XbG_H273<=Vw;
XbG_H274<=Vw;
XbG_H275<=Vw;
XbG_H276<=Vw;
XbG_H277<=Vw;
XbG_H278<=Vw;
XbG_H279<=Vw;
XbG_H28<=Vw;
XbG_H280<=Vw;
XbG_H281<=Vw;
XbG_H282<=Vw;
XbG_H283<=Vw;
XbG_H284<=Vw;
XbG_H285<=Vw;
XbG_H286<=Vw;
XbG_H287<=Vw;
XbG_H288<=Vw;
XbG_H289<=Vw;
XbG_H29<=Vw;
XbG_H290<=Vw;
XbG_H291<=Vw;
XbG_H292<=Vw;
XbG_H293<=Vw;
XbG_H294<=Vw;
XbG_H295<=Vw;
XbG_H296<=Vw;
XbG_H297<=Vw;
XbG_H298<=Vw;
XbG_H299<=Vw;
XbG_H3<=Vw;
XbG_H30<=Vw;
XbG_H300<=Vw;
XbG_H301<=Vw;
XbG_H302<=Vw;
XbG_H303<=Vw;
XbG_H304<=Vw;
XbG_H305<=Vw;
XbG_H306<=Vw;
XbG_H307<=Vw;
XbG_H308<=Vw;
XbG_H309<=Vw;
XbG_H31<=Vw;
XbG_H310<=Vw;
XbG_H311<=Vw;
XbG_H312<=Vw;
XbG_H313<=Vw;
XbG_H314<=Vw;
XbG_H315<=Vw;
XbG_H316<=Vw;
XbG_H317<=Vw;
XbG_H318<=Vw;
XbG_H319<=Vw;
XbG_H32<=Vw;
XbG_H320<=Vw;
XbG_H321<=Vw;
XbG_H322<=Vw;
XbG_H323<=Vw;
XbG_H324<=Vw;
XbG_H325<=Vw;
XbG_H326<=Vw;
XbG_H327<=Vw;
XbG_H328<=Vw;
XbG_H329<=Vw;
XbG_H33<=Vw;
XbG_H330<=Vw;
XbG_H331<=Vw;
XbG_H332<=Vw;
XbG_H333<=Vw;
XbG_H334<=Vw;
XbG_H335<=Vw;
XbG_H336<=Vw;
XbG_H337<=Vw;
XbG_H338<=Vw;
XbG_H339<=Vw;
XbG_H34<=Vw;
XbG_H340<=Vw;
XbG_H341<=Vw;
XbG_H342<=Vw;
XbG_H343<=Vw;
XbG_H344<=Vw;
XbG_H345<=Vw;
XbG_H346<=Vw;
XbG_H347<=Vw;
XbG_H348<=Vw;
XbG_H349<=Vw;
XbG_H35<=Vw;
XbG_H350<=Vw;
XbG_H351<=Vw;
XbG_H352<=Vw;
XbG_H353<=Vw;
XbG_H354<=Vw;
XbG_H355<=Vw;
XbG_H356<=Vw;
XbG_H357<=Vw;
XbG_H358<=Vw;
XbG_H359<=Vw;
XbG_H36<=Vw;
XbG_H360<=Vw;
XbG_H361<=Vw;
XbG_H362<=Vw;
XbG_H363<=Vw;
XbG_H364<=Vw;
XbG_H365<=Vw;
XbG_H366<=Vw;
XbG_H367<=Vw;
XbG_H368<=Vw;
XbG_H369<=Vw;
XbG_H37<=Vw;
XbG_H370<=Vw;
XbG_H371<=Vw;
XbG_H372<=Vw;
XbG_H373<=Vw;
XbG_H374<=Vw;
XbG_H375<=Vw;
XbG_H376<=Vw;
XbG_H377<=Vw;
XbG_H378<=Vw;
XbG_H379<=Vw;
XbG_H38<=Vw;
XbG_H380<=Vw;
XbG_H381<=Vw;
XbG_H382<=Vw;
XbG_H383<=Vw;
XbG_H384<=Vw;
XbG_H385<=Vw;
XbG_H386<=Vw;
XbG_H387<=Vw;
XbG_H388<=Vw;
XbG_H389<=Vw;
XbG_H39<=Vw;
XbG_H390<=Vw;
XbG_H391<=Vw;
XbG_H392<=Vw;
XbG_H393<=Vw;
XbG_H394<=Vw;
XbG_H395<=Vw;
XbG_H396<=Vw;
XbG_H397<=Vw;
XbG_H398<=Vw;
XbG_H399<=Vw;
XbG_H4<=Vw;
XbG_H40<=Vw;
XbG_H400<=Vw;
XbG_H401<=Vw;
XbG_H402<=Vw;
XbG_H403<=Vw;
XbG_H404<=Vw;
XbG_H405<=Vw;
XbG_H406<=Vw;
XbG_H407<=Vw;
XbG_H408<=Vw;
XbG_H409<=Vw;
XbG_H41<=Vw;
XbG_H410<=Vw;
XbG_H411<=Vw;
XbG_H412<=Vw;
XbG_H413<=Vw;
XbG_H414<=Vw;
XbG_H415<=Vw;
XbG_H416<=Vw;
XbG_H417<=Vw;
XbG_H418<=Vw;
XbG_H419<=Vw;
XbG_H42<=Vw;
XbG_H420<=Vw;
XbG_H421<=Vw;
XbG_H422<=Vw;
XbG_H423<=Vw;
XbG_H424<=Vw;
XbG_H425<=Vw;
XbG_H426<=Vw;
XbG_H427<=Vw;
XbG_H428<=Vw;
XbG_H429<=Vw;
XbG_H43<=Vw;
XbG_H430<=Vw;
XbG_H431<=Vw;
XbG_H432<=Vw;
XbG_H433<=Vw;
XbG_H434<=Vw;
XbG_H435<=Vw;
XbG_H436<=Vw;
XbG_H437<=Vw;
XbG_H438<=Vw;
XbG_H439<=Vw;
XbG_H44<=Vw;
XbG_H440<=Vw;
XbG_H441<=Vw;
XbG_H442<=Vw;
XbG_H443<=Vw;
XbG_H444<=Vw;
XbG_H445<=Vw;
XbG_H446<=Vw;
XbG_H447<=Vw;
XbG_H448<=Vw;
XbG_H449<=Vw;
XbG_H45<=Vw;
XbG_H450<=Vw;
XbG_H451<=Vw;
XbG_H452<=Vw;
XbG_H453<=Vw;
XbG_H454<=Vw;
XbG_H455<=Vw;
XbG_H456<=Vw;
XbG_H457<=Vw;
XbG_H458<=Vw;
XbG_H459<=Vw;
XbG_H46<=Vw;
XbG_H460<=Vw;
XbG_H461<=Vw;
XbG_H462<=Vw;
XbG_H463<=Vw;
XbG_H464<=Vw;
XbG_H465<=Vw;
XbG_H466<=Vw;
XbG_H467<=Vw;
XbG_H468<=Vw;
XbG_H469<=Vw;
XbG_H47<=Vw;
XbG_H470<=Vw;
XbG_H471<=Vw;
XbG_H472<=Vw;
XbG_H473<=Vw;
XbG_H474<=Vw;
XbG_H475<=Vw;
XbG_H476<=Vw;
XbG_H477<=Vw;
XbG_H478<=Vw;
XbG_H479<=Vw;
XbG_H48<=Vw;
XbG_H480<=Vw;
XbG_H481<=Vw;
XbG_H482<=Vw;
XbG_H483<=Vw;
XbG_H484<=Vw;
XbG_H485<=Vw;
XbG_H486<=Vw;
XbG_H487<=Vw;
XbG_H488<=Vw;
XbG_H489<=Vw;
XbG_H49<=Vw;
XbG_H490<=Vw;
XbG_H491<=Vw;
XbG_H492<=Vw;
XbG_H493<=Vw;
XbG_H494<=Vw;
XbG_H495<=Vw;
XbG_H496<=Vw;
XbG_H497<=Vw;
XbG_H498<=Vw;
XbG_H499<=Vw;
XbG_H5<=Vw;
XbG_H50<=Vw;
XbG_H500<=Vw;
XbG_H501<=Vw;
XbG_H502<=Vw;
XbG_H503<=Vw;
XbG_H504<=Vw;
XbG_H505<=Vw;
XbG_H506<=Vw;
XbG_H507<=Vw;
XbG_H508<=Vw;
XbG_H509<=Vw;
XbG_H51<=Vw;
XbG_H510<=Vw;
XbG_H511<=Vw;
XbG_H512<=Vw;
XbG_H513<=Vw;
XbG_H514<=Vw;
XbG_H515<=Vw;
XbG_H516<=Vw;
XbG_H517<=Vw;
XbG_H518<=Vw;
XbG_H519<=Vw;
XbG_H52<=Vw;
XbG_H520<=Vw;
XbG_H521<=Vw;
XbG_H522<=Vw;
XbG_H523<=Vw;
XbG_H524<=Vw;
XbG_H525<=Vw;
XbG_H526<=Vw;
XbG_H527<=Vw;
XbG_H528<=Vw;
XbG_H529<=Vw;
XbG_H53<=Vw;
XbG_H530<=Vw;
XbG_H531<=Vw;
XbG_H532<=Vw;
XbG_H533<=Vw;
XbG_H534<=Vw;
XbG_H535<=Vw;
XbG_H536<=Vw;
XbG_H537<=Vw;
XbG_H538<=Vw;
XbG_H539<=Vw;
XbG_H54<=Vw;
XbG_H540<=Vw;
XbG_H541<=Vw;
XbG_H542<=Vw;
XbG_H543<=Vw;
XbG_H544<=Vw;
XbG_H545<=Vw;
XbG_H546<=Vw;
XbG_H547<=Vw;
XbG_H548<=Vw;
XbG_H549<=Vw;
XbG_H55<=Vw;
XbG_H550<=Vw;
XbG_H551<=Vw;
XbG_H552<=Vw;
XbG_H553<=Vw;
XbG_H554<=Vw;
XbG_H555<=Vw;
XbG_H556<=Vw;
XbG_H557<=Vw;
XbG_H558<=Vw;
XbG_H559<=Vw;
XbG_H56<=Vw;
XbG_H560<=Vw;
XbG_H561<=Vw;
XbG_H562<=Vw;
XbG_H563<=Vw;
XbG_H564<=Vw;
XbG_H565<=Vw;
XbG_H566<=Vw;
XbG_H567<=Vw;
XbG_H568<=Vw;
XbG_H569<=Vw;
XbG_H57<=Vw;
XbG_H570<=Vw;
XbG_H571<=Vw;
XbG_H572<=Vw;
XbG_H573<=Vw;
XbG_H574<=Vw;
XbG_H575<=Vw;
XbG_H576<=Vw;
XbG_H577<=Vw;
XbG_H578<=Vw;
XbG_H579<=Vw;
XbG_H58<=Vw;
XbG_H580<=Vw;
XbG_H581<=Vw;
XbG_H582<=Vw;
XbG_H583<=Vw;
XbG_H584<=Vw;
XbG_H585<=Vw;
XbG_H586<=Vw;
XbG_H587<=Vw;
XbG_H588<=Vw;
XbG_H589<=Vw;
XbG_H59<=Vw;
XbG_H590<=Vw;
XbG_H591<=Vw;
XbG_H592<=Vw;
XbG_H593<=Vw;
XbG_H594<=Vw;
XbG_H595<=Vw;
XbG_H596<=Vw;
XbG_H597<=Vw;
XbG_H598<=Vw;
XbG_H599<=Vw;
XbG_H6<=Vw;
XbG_H60<=Vw;
XbG_H600<=Vw;
XbG_H601<=Vw;
XbG_H602<=Vw;
XbG_H603<=Vw;
XbG_H604<=Vw;
XbG_H605<=Vw;
XbG_H606<=Vw;
XbG_H607<=Vw;
XbG_H608<=Vw;
XbG_H609<=Vw;
XbG_H61<=Vw;
XbG_H610<=Vw;
XbG_H611<=Vw;
XbG_H612<=Vw;
XbG_H613<=Vw;
XbG_H614<=Vw;
XbG_H615<=Vw;
XbG_H616<=Vw;
XbG_H617<=Vw;
XbG_H618<=Vw;
XbG_H619<=Vw;
XbG_H62<=Vw;
XbG_H620<=Vw;
XbG_H621<=Vw;
XbG_H622<=Vw;
XbG_H623<=Vw;
XbG_H624<=Vw;
XbG_H625<=Vw;
XbG_H626<=Vw;
XbG_H627<=Vw;
XbG_H628<=Vw;
XbG_H629<=Vw;
XbG_H63<=Vw;
XbG_H630<=Vw;
XbG_H631<=Vw;
XbG_H632<=Vw;
XbG_H633<=Vw;
XbG_H634<=Vw;
XbG_H635<=Vw;
XbG_H636<=Vw;
XbG_H637<=Vw;
XbG_H638<=Vw;
XbG_H639<=Vw;
XbG_H64<=Vw;
XbG_H640<=Vw;
XbG_H641<=Vw;
XbG_H642<=Vw;
XbG_H643<=Vw;
XbG_H644<=Vw;
XbG_H645<=Vw;
XbG_H646<=Vw;
XbG_H647<=Vw;
XbG_H648<=Vw;
XbG_H649<=Vw;
XbG_H65<=Vw;
XbG_H650<=Vw;
XbG_H651<=Vw;
XbG_H652<=Vw;
XbG_H653<=Vw;
XbG_H654<=Vw;
XbG_H655<=Vw;
XbG_H656<=Vw;
XbG_H657<=Vw;
XbG_H658<=Vw;
XbG_H659<=Vw;
XbG_H66<=Vw;
XbG_H660<=Vw;
XbG_H661<=zero;
XbG_H662<=zero;
XbG_H663<=zero;
XbG_H664<=zero;
XbG_H665<=zero;
XbG_H666<=zero;
XbG_H667<=zero;
XbG_H668<=zero;
XbG_H669<=zero;
XbG_H67<=Vw;
XbG_H670<=zero;
XbG_H671<=zero;
XbG_H672<=zero;
XbG_H673<=zero;
XbG_H674<=zero;
XbG_H675<=zero;
XbG_H676<=zero;
XbG_H677<=zero;
XbG_H678<=zero;
XbG_H679<=zero;
XbG_H68<=Vw;
XbG_H680<=zero;
XbG_H681<=zero;
XbG_H682<=zero;
XbG_H683<=zero;
XbG_H684<=zero;
XbG_H685<=zero;
XbG_H686<=zero;
XbG_H687<=zero;
XbG_H688<=zero;
XbG_H689<=zero;
XbG_H69<=Vw;
XbG_H690<=zero;
XbG_H691<=zero;
XbG_H692<=zero;
XbG_H693<=zero;
XbG_H694<=zero;
XbG_H695<=zero;
XbG_H696<=zero;
XbG_H697<=zero;
XbG_H698<=zero;
XbG_H699<=zero;
XbG_H7<=Vw;
XbG_H70<=Vw;
XbG_H700<=zero;
XbG_H701<=zero;
XbG_H702<=zero;
XbG_H703<=zero;
XbG_H704<=zero;
XbG_H705<=zero;
XbG_H706<=zero;
XbG_H707<=zero;
XbG_H708<=zero;
XbG_H709<=zero;
XbG_H71<=Vw;
XbG_H710<=zero;
XbG_H711<=zero;
XbG_H712<=zero;
XbG_H713<=zero;
XbG_H714<=zero;
XbG_H715<=zero;
XbG_H716<=zero;
XbG_H717<=zero;
XbG_H718<=zero;
XbG_H719<=zero;
XbG_H72<=Vw;
XbG_H720<=zero;
XbG_H721<=zero;
XbG_H722<=Vw;
XbG_H723<=Vw;
XbG_H724<=Vw;
XbG_H725<=Vw;
XbG_H726<=Vw;
XbG_H727<=Vw;
XbG_H728<=Vw;
XbG_H729<=Vw;
XbG_H73<=Vw;
XbG_H730<=Vw;
XbG_H731<=Vw;
XbG_H732<=Vw;
XbG_H733<=Vw;
XbG_H734<=Vw;
XbG_H735<=Vw;
XbG_H74<=Vw;
XbG_H75<=Vw;
XbG_H76<=Vw;
XbG_H77<=Vw;
XbG_H78<=Vw;
XbG_H79<=Vw;
XbG_H8<=Vw;
XbG_H80<=Vw;
XbG_H81<=Vw;
XbG_H82<=Vw;
XbG_H83<=Vw;
XbG_H84<=Vw;
XbG_H85<=Vw;
XbG_H86<=Vw;
XbG_H87<=Vw;
XbG_H88<=Vw;
XbG_H89<=Vw;
XbG_H9<=Vw;
XbG_H90<=Vw;
XbG_H91<=Vw;
XbG_H92<=Vw;
XbG_H93<=Vw;
XbG_H94<=Vw;
XbG_H95<=Vw;
XbG_H96<=Vw;
XbG_H97<=Vw;
XbG_H98<=Vw;
XbG_H99<=Vw;
XbG_V0<=zero;
XbG_V1<=zero;
XbG_V10<=zero;
XbG_V100<=Vr;
XbG_V101<=Vr, (others=>'Z') after 1 ps;
XbG_V102<=Vr;
XbG_V103<=Vr, (others=>'Z') after 1 ps;
XbG_V104<=Vr;
XbG_V105<=Vr, (others=>'Z') after 1 ps;
XbG_V106<=Vr;
XbG_V107<=Vr, (others=>'Z') after 1 ps;
XbG_V108<=Vr;
XbG_V109<=Vr, (others=>'Z') after 1 ps;
XbG_V11<=zero;
XbG_V110<=Vr;
XbG_V111<=Vr, (others=>'Z') after 1 ps;
XbG_V112<=Vr;
XbG_V113<=Vr, (others=>'Z') after 1 ps;
XbG_V114<=Vr;
XbG_V115<=Vr, (others=>'Z') after 1 ps;
XbG_V116<=Vr;
XbG_V117<=Vr, (others=>'Z') after 1 ps;
XbG_V118<=Vr;
XbG_V119<=Vr, (others=>'Z') after 1 ps;
XbG_V12<=zero;
XbG_V120<=Vr;
XbG_V121<=Vr, (others=>'Z') after 1 ps;
XbG_V122<=Vr;
XbG_V123<=Vr, (others=>'Z') after 1 ps;
XbG_V124<=Vr;
XbG_V125<=Vr, (others=>'Z') after 1 ps;
XbG_V126<=Vr;
XbG_V127<=Vr, (others=>'Z') after 1 ps;
XbG_V128<=Vr;
XbG_V129<=Vr, (others=>'Z') after 1 ps;
XbG_V13<=zero;
XbG_V130<=Vr;
XbG_V131<=Vr, (others=>'Z') after 1 ps;
XbG_V132<=Vr;
XbG_V133<=Vr, (others=>'Z') after 1 ps;
XbG_V134<=Vr;
XbG_V135<=Vr, (others=>'Z') after 1 ps;
XbG_V136<=Vr;
XbG_V137<=Vr, (others=>'Z') after 1 ps;
XbG_V138<=Vr;
XbG_V139<=Vr, (others=>'Z') after 1 ps;
XbG_V14<=zero;
XbG_V140<=Vr;
XbG_V141<=Vr, (others=>'Z') after 1 ps;
XbG_V142<=Vr;
XbG_V143<=Vr, (others=>'Z') after 1 ps;
XbG_V144<=Vr;
XbG_V145<=Vr, (others=>'Z') after 1 ps;
XbG_V146<=Vr;
XbG_V147<=Vr, (others=>'Z') after 1 ps;
XbG_V148<=Vr;
XbG_V149<=Vr, (others=>'Z') after 1 ps;
XbG_V15<=zero;
XbG_V150<=Vr;
XbG_V151<=Vr, (others=>'Z') after 1 ps;
XbG_V152<=Vr;
XbG_V153<=Vr, (others=>'Z') after 1 ps;
XbG_V154<=Vr;
XbG_V155<=Vr, (others=>'Z') after 1 ps;
XbG_V156<=Vr;
XbG_V157<=Vr, (others=>'Z') after 1 ps;
XbG_V158<=Vr;
XbG_V159<=Vr, (others=>'Z') after 1 ps;
XbG_V16<=zero;
XbG_V160<=Vr;
XbG_V161<=Vr, (others=>'Z') after 1 ps;
XbG_V162<=Vr;
XbG_V163<=Vr, (others=>'Z') after 1 ps;
XbG_V164<=Vr;
XbG_V165<=Vr, (others=>'Z') after 1 ps;
XbG_V166<=Vr;
XbG_V167<=Vr, (others=>'Z') after 1 ps;
XbG_V168<=Vr;
XbG_V169<=Vr, (others=>'Z') after 1 ps;
XbG_V17<=zero;
XbG_V170<=Vr;
XbG_V171<=Vr, (others=>'Z') after 1 ps;
XbG_V172<=Vr;
XbG_V173<=Vr, (others=>'Z') after 1 ps;
XbG_V174<=Vr;
XbG_V175<=Vr, (others=>'Z') after 1 ps;
XbG_V176<=Vr;
XbG_V177<=Vr, (others=>'Z') after 1 ps;
XbG_V178<=Vr;
XbG_V179<=Vr, (others=>'Z') after 1 ps;
XbG_V18<=zero;
XbG_V180<=Vr;
XbG_V181<=Vr, (others=>'Z') after 1 ps;
XbG_V182<=Vr;
XbG_V183<=Vr, (others=>'Z') after 1 ps;
XbG_V184<=Vr;
XbG_V185<=Vr, (others=>'Z') after 1 ps;
XbG_V186<=Vr;
XbG_V187<=Vr, (others=>'Z') after 1 ps;
XbG_V188<=Vr;
XbG_V189<=Vr, (others=>'Z') after 1 ps;
XbG_V19<=zero;
XbG_V2<=zero;
XbG_V20<=zero;
XbG_V21<=zero;
XbG_V22<=zero;
XbG_V23<=zero;
XbG_V24<=zero;
XbG_V25<=zero;
XbG_V26<=zero;
XbG_V27<=zero;
XbG_V28<=zero;
XbG_V29<=zero;
XbG_V3<=zero;
XbG_V30<=zero;
XbG_V31<=zero;
XbG_V32<=zero;
XbG_V33<=zero;
XbG_V34<=zero;
XbG_V35<=zero;
XbG_V36<=zero;
XbG_V37<=zero;
XbG_V38<=zero;
XbG_V39<=zero;
XbG_V4<=zero;
XbG_V40<=zero;
XbG_V41<=zero;
XbG_V42<=zero;
XbG_V43<=zero;
XbG_V44<=zero;
XbG_V45<=zero;
XbG_V46<=zero;
XbG_V47<=zero;
XbG_V48<=zero;
XbG_V49<=zero;
XbG_V5<=zero;
XbG_V50<=zero;
XbG_V51<=zero;
XbG_V52<=zero;
XbG_V53<=zero;
XbG_V54<=zero;
XbG_V55<=zero;
XbG_V56<=zero;
XbG_V57<=zero;
XbG_V58<=zero;
XbG_V59<=zero;
XbG_V6<=zero;
XbG_V60<=zero;
XbG_V61<=zero;
XbG_V62<=zero;
XbG_V63<=zero;
XbG_V64<=zero;
XbG_V65<=zero;
XbG_V66<=zero;
XbG_V67<=zero;
XbG_V68<=Vr;
XbG_V69<=Vr, (others=>'Z') after 1 ps;
XbG_V7<=zero;
XbG_V70<=Vr;
XbG_V71<=Vr, (others=>'Z') after 1 ps;
XbG_V72<=Vr;
XbG_V73<=Vr, (others=>'Z') after 1 ps;
XbG_V74<=Vr;
XbG_V75<=Vr, (others=>'Z') after 1 ps;
XbG_V76<=Vr;
XbG_V77<=Vr, (others=>'Z') after 1 ps;
XbG_V78<=Vr;
XbG_V79<=Vr, (others=>'Z') after 1 ps;
XbG_V8<=zero;
XbG_V80<=Vr;
XbG_V81<=Vr, (others=>'Z') after 1 ps;
XbG_V82<=Vr;
XbG_V83<=Vr, (others=>'Z') after 1 ps;
XbG_V84<=Vr;
XbG_V85<=Vr, (others=>'Z') after 1 ps;
XbG_V86<=Vr;
XbG_V87<=Vr, (others=>'Z') after 1 ps;
XbG_V88<=Vr;
XbG_V89<=Vr, (others=>'Z') after 1 ps;
XbG_V9<=zero;
XbG_V90<=Vr;
XbG_V91<=Vr, (others=>'Z') after 1 ps;
XbG_V92<=Vr;
XbG_V93<=Vr, (others=>'Z') after 1 ps;
XbG_V94<=Vr;
XbG_V95<=Vr, (others=>'Z') after 1 ps;
XbG_V96<=Vr;
XbG_V97<=Vr, (others=>'Z') after 1 ps;
XbG_V98<=Vr;
XbG_V99<=Vr, (others=>'Z') after 1 ps;

next_state<=F_INR;

when F_INR =>

XbG_H0<=Vr;
XbG_H1<=Vr;
XbG_H10<=Vr;
XbG_H100<=Vr;
XbG_H101<=Vr;
XbG_H102<=Vr;
XbG_H103<=Vr;
XbG_H104<=Vr;
XbG_H105<=Vr;
XbG_H106<=Vr;
XbG_H107<=Vr;
XbG_H108<=Vr;
XbG_H109<=Vr;
XbG_H11<=Vr;
XbG_H110<=Vr;
XbG_H111<=Vr;
XbG_H112<=Vr;
XbG_H113<=Vr;
XbG_H114<=Vr;
XbG_H115<=Vr;
XbG_H116<=Vr;
XbG_H117<=Vr;
XbG_H118<=Vr;
XbG_H119<=Vr;
XbG_H12<=Vr;
XbG_H120<=Vr;
XbG_H121<=Vr;
XbG_H122<=Vr;
XbG_H123<=Vr;
XbG_H124<=Vr;
XbG_H125<=Vr;
XbG_H126<=Vr;
XbG_H127<=Vr;
XbG_H128<=Vr;
XbG_H129<=Vr;
XbG_H13<=Vr;
XbG_H130<=Vr;
XbG_H131<=Vr;
XbG_H132<=Vr;
XbG_H133<=Vr;
XbG_H134<=Vr;
XbG_H135<=Vr;
XbG_H136<=Vr;
XbG_H137<=Vr;
XbG_H138<=Vr;
XbG_H139<=Vr;
XbG_H14<=Vr;
XbG_H140<=Vr;
XbG_H141<=Vr;
XbG_H142<=Vr;
XbG_H143<=Vr;
XbG_H144<=Vr;
XbG_H145<=Vr;
XbG_H146<=Vr;
XbG_H147<=Vr;
XbG_H148<=Vr;
XbG_H149<=Vr;
XbG_H15<=Vr;
XbG_H150<=Vr;
XbG_H151<=Vr;
XbG_H152<=Vr;
XbG_H153<=Vr;
XbG_H154<=Vr;
XbG_H155<=Vr;
XbG_H156<=Vr;
XbG_H157<=Vr;
XbG_H158<=Vr;
XbG_H159<=Vr;
XbG_H16<=Vr;
XbG_H160<=Vr;
XbG_H161<=Vr;
XbG_H162<=Vr;
XbG_H163<=Vr;
XbG_H164<=Vr;
XbG_H165<=Vr;
XbG_H166<=Vr;
XbG_H167<=Vr;
XbG_H168<=Vr;
XbG_H169<=Vr;
XbG_H17<=Vr;
XbG_H170<=Vr;
XbG_H171<=Vr;
XbG_H172<=Vr;
XbG_H173<=Vr;
XbG_H174<=Vr;
XbG_H175<=Vr;
XbG_H176<=Vr;
XbG_H177<=Vr;
XbG_H178<=Vr;
XbG_H179<=Vr;
XbG_H18<=Vr;
XbG_H180<=Vr;
XbG_H181<=Vr;
XbG_H182<=Vr;
XbG_H183<=Vr;
XbG_H184<=Vr;
XbG_H185<=Vr;
XbG_H186<=Vr;
XbG_H187<=Vr;
XbG_H188<=Vr;
XbG_H189<=Vr;
XbG_H19<=Vr;
XbG_H190<=Vr;
XbG_H191<=Vr;
XbG_H192<=Vr;
XbG_H193<=Vr;
XbG_H194<=Vr;
XbG_H195<=Vr;
XbG_H196<=Vr;
XbG_H197<=Vr;
XbG_H198<=Vr;
XbG_H199<=Vr;
XbG_H2<=Vr;
XbG_H20<=Vr;
XbG_H200<=Vr;
XbG_H201<=Vr;
XbG_H202<=Vr;
XbG_H203<=Vr;
XbG_H204<=Vr;
XbG_H205<=Vr;
XbG_H206<=Vr;
XbG_H207<=Vr;
XbG_H208<=Vr;
XbG_H209<=Vr;
XbG_H21<=Vr;
XbG_H210<=Vr;
XbG_H211<=Vr;
XbG_H212<=Vr;
XbG_H213<=Vr;
XbG_H214<=Vr;
XbG_H215<=Vr;
XbG_H216<=Vr;
XbG_H217<=Vr;
XbG_H218<=Vr;
XbG_H219<=Vr;
XbG_H22<=Vr;
XbG_H220<=Vr;
XbG_H221<=Vr;
XbG_H222<=Vr;
XbG_H223<=Vr;
XbG_H224<=Vr;
XbG_H225<=Vr;
XbG_H226<=Vr;
XbG_H227<=Vr;
XbG_H228<=Vr;
XbG_H229<=Vr;
XbG_H23<=Vr;
XbG_H230<=Vr;
XbG_H231<=Vr;
XbG_H232<=Vr;
XbG_H233<=Vr;
XbG_H234<=Vr;
XbG_H235<=Vr;
XbG_H236<=Vr;
XbG_H237<=Vr;
XbG_H238<=Vr;
XbG_H239<=Vr;
XbG_H24<=Vr;
XbG_H240<=Vr;
XbG_H241<=Vr;
XbG_H242<=Vr;
XbG_H243<=Vr;
XbG_H244<=Vr;
XbG_H245<=Vr;
XbG_H246<=Vr;
XbG_H247<=Vr;
XbG_H248<=Vr;
XbG_H249<=Vr;
XbG_H25<=Vr;
XbG_H250<=Vr;
XbG_H251<=Vr;
XbG_H252<=Vr;
XbG_H253<=Vr;
XbG_H254<=Vr;
XbG_H255<=Vr;
XbG_H256<=Vr;
XbG_H257<=Vr;
XbG_H258<=Vr;
XbG_H259<=Vr;
XbG_H26<=Vr;
XbG_H260<=Vr;
XbG_H261<=Vr;
XbG_H262<=Vr;
XbG_H263<=Vr;
XbG_H264<=Vr;
XbG_H265<=Vr;
XbG_H266<=Vr;
XbG_H267<=Vr;
XbG_H268<=Vr;
XbG_H269<=Vr;
XbG_H27<=Vr;
XbG_H270<=Vr;
XbG_H271<=Vr;
XbG_H272<=Vr;
XbG_H273<=Vr;
XbG_H274<=Vr;
XbG_H275<=Vr;
XbG_H276<=Vr;
XbG_H277<=Vr;
XbG_H278<=Vr;
XbG_H279<=Vr;
XbG_H28<=Vr;
XbG_H280<=Vr;
XbG_H281<=Vr;
XbG_H282<=Vr;
XbG_H283<=Vr;
XbG_H284<=Vr;
XbG_H285<=Vr;
XbG_H286<=Vr;
XbG_H287<=Vr;
XbG_H288<=Vr;
XbG_H289<=Vr;
XbG_H29<=Vr;
XbG_H290<=Vr;
XbG_H291<=Vr;
XbG_H292<=Vr;
XbG_H293<=Vr;
XbG_H294<=Vr;
XbG_H295<=Vr;
XbG_H296<=Vr;
XbG_H297<=Vr;
XbG_H298<=Vr;
XbG_H299<=Vr;
XbG_H3<=Vr;
XbG_H30<=Vr;
XbG_H300<=Vr;
XbG_H301<=Vr;
XbG_H302<=Vr;
XbG_H303<=Vr;
XbG_H304<=Vr;
XbG_H305<=Vr;
XbG_H306<=Vr;
XbG_H307<=Vr;
XbG_H308<=Vr;
XbG_H309<=Vr;
XbG_H31<=Vr;
XbG_H310<=Vr;
XbG_H311<=Vr;
XbG_H312<=Vr;
XbG_H313<=Vr;
XbG_H314<=Vr;
XbG_H315<=Vr;
XbG_H316<=Vr;
XbG_H317<=Vr;
XbG_H318<=Vr;
XbG_H319<=Vr;
XbG_H32<=Vr;
XbG_H320<=Vr;
XbG_H321<=Vr;
XbG_H322<=Vr;
XbG_H323<=Vr;
XbG_H324<=Vr;
XbG_H325<=Vr;
XbG_H326<=Vr;
XbG_H327<=Vr;
XbG_H328<=Vr;
XbG_H329<=Vr;
XbG_H33<=Vr;
XbG_H330<=Vr;
XbG_H331<=Vr;
XbG_H332<=Vr;
XbG_H333<=Vr;
XbG_H334<=Vr;
XbG_H335<=Vr;
XbG_H336<=Vr;
XbG_H337<=Vr;
XbG_H338<=Vr;
XbG_H339<=Vr;
XbG_H34<=Vr;
XbG_H340<=Vr;
XbG_H341<=Vr;
XbG_H342<=Vr;
XbG_H343<=Vr;
XbG_H344<=Vr;
XbG_H345<=Vr;
XbG_H346<=Vr;
XbG_H347<=Vr;
XbG_H348<=Vr;
XbG_H349<=Vr;
XbG_H35<=Vr;
XbG_H350<=Vr;
XbG_H351<=Vr;
XbG_H352<=Vr;
XbG_H353<=Vr;
XbG_H354<=Vr;
XbG_H355<=Vr;
XbG_H356<=Vr;
XbG_H357<=Vr;
XbG_H358<=Vr;
XbG_H359<=Vr;
XbG_H36<=Vr;
XbG_H360<=Vr;
XbG_H361<=Vr;
XbG_H362<=Vr;
XbG_H363<=Vr;
XbG_H364<=Vr;
XbG_H365<=Vr;
XbG_H366<=Vr;
XbG_H367<=Vr;
XbG_H368<=Vr;
XbG_H369<=Vr;
XbG_H37<=Vr;
XbG_H370<=Vr;
XbG_H371<=Vr;
XbG_H372<=Vr;
XbG_H373<=Vr;
XbG_H374<=Vr;
XbG_H375<=Vr;
XbG_H376<=Vr;
XbG_H377<=Vr;
XbG_H378<=Vr;
XbG_H379<=Vr;
XbG_H38<=Vr;
XbG_H380<=Vr;
XbG_H381<=Vr;
XbG_H382<=Vr;
XbG_H383<=Vr;
XbG_H384<=Vr;
XbG_H385<=Vr;
XbG_H386<=Vr;
XbG_H387<=Vr;
XbG_H388<=Vr;
XbG_H389<=Vr;
XbG_H39<=Vr;
XbG_H390<=Vr;
XbG_H391<=Vr;
XbG_H392<=Vr;
XbG_H393<=Vr;
XbG_H394<=Vr;
XbG_H395<=Vr;
XbG_H396<=Vr;
XbG_H397<=Vr;
XbG_H398<=Vr;
XbG_H399<=Vr;
XbG_H4<=Vr;
XbG_H40<=Vr;
XbG_H400<=Vr;
XbG_H401<=Vr;
XbG_H402<=Vr;
XbG_H403<=Vr;
XbG_H404<=Vr;
XbG_H405<=Vr;
XbG_H406<=Vr;
XbG_H407<=Vr;
XbG_H408<=Vr;
XbG_H409<=Vr;
XbG_H41<=Vr;
XbG_H410<=Vr;
XbG_H411<=Vr;
XbG_H412<=Vr;
XbG_H413<=Vr;
XbG_H414<=Vr;
XbG_H415<=Vr;
XbG_H416<=Vr;
XbG_H417<=Vr;
XbG_H418<=Vr;
XbG_H419<=Vr;
XbG_H42<=Vr;
XbG_H420<=Vr;
XbG_H421<=Vr;
XbG_H422<=Vr;
XbG_H423<=Vr;
XbG_H424<=Vr;
XbG_H425<=Vr;
XbG_H426<=Vr;
XbG_H427<=Vr;
XbG_H428<=Vr;
XbG_H429<=Vr;
XbG_H43<=Vr;
XbG_H430<=Vr;
XbG_H431<=Vr;
XbG_H432<=Vr;
XbG_H433<=Vr;
XbG_H434<=Vr;
XbG_H435<=Vr;
XbG_H436<=Vr;
XbG_H437<=Vr;
XbG_H438<=Vr;
XbG_H439<=Vr;
XbG_H44<=Vr;
XbG_H440<=Vr;
XbG_H441<=Vr;
XbG_H442<=Vr;
XbG_H443<=Vr;
XbG_H444<=Vr;
XbG_H445<=Vr;
XbG_H446<=Vr;
XbG_H447<=Vr;
XbG_H448<=Vr;
XbG_H449<=Vr;
XbG_H45<=Vr;
XbG_H450<=Vr;
XbG_H451<=Vr;
XbG_H452<=Vr;
XbG_H453<=Vr;
XbG_H454<=Vr;
XbG_H455<=Vr;
XbG_H456<=Vr;
XbG_H457<=Vr;
XbG_H458<=Vr;
XbG_H459<=Vr;
XbG_H46<=Vr;
XbG_H460<=Vr;
XbG_H461<=Vr;
XbG_H462<=Vr;
XbG_H463<=Vr;
XbG_H464<=Vr;
XbG_H465<=Vr;
XbG_H466<=Vr;
XbG_H467<=Vr;
XbG_H468<=Vr;
XbG_H469<=Vr;
XbG_H47<=Vr;
XbG_H470<=Vr;
XbG_H471<=Vr;
XbG_H472<=Vr;
XbG_H473<=Vr;
XbG_H474<=Vr;
XbG_H475<=Vr;
XbG_H476<=Vr;
XbG_H477<=Vr;
XbG_H478<=Vr;
XbG_H479<=Vr;
XbG_H48<=Vr;
XbG_H480<=Vr;
XbG_H481<=Vr;
XbG_H482<=Vr;
XbG_H483<=Vr;
XbG_H484<=Vr;
XbG_H485<=Vr;
XbG_H486<=Vr;
XbG_H487<=Vr;
XbG_H488<=Vr;
XbG_H489<=Vr;
XbG_H49<=Vr;
XbG_H490<=Vr;
XbG_H491<=Vr;
XbG_H492<=Vr;
XbG_H493<=Vr;
XbG_H494<=Vr;
XbG_H495<=Vr;
XbG_H496<=Vr;
XbG_H497<=Vr;
XbG_H498<=Vr;
XbG_H499<=Vr;
XbG_H5<=Vr;
XbG_H50<=Vr;
XbG_H500<=Vr;
XbG_H501<=Vr;
XbG_H502<=Vr;
XbG_H503<=Vr;
XbG_H504<=Vr;
XbG_H505<=Vr;
XbG_H506<=Vr;
XbG_H507<=Vr;
XbG_H508<=Vr;
XbG_H509<=Vr;
XbG_H51<=Vr;
XbG_H510<=Vr;
XbG_H511<=Vr;
XbG_H512<=Vr;
XbG_H513<=Vr;
XbG_H514<=Vr;
XbG_H515<=Vr;
XbG_H516<=Vr;
XbG_H517<=Vr;
XbG_H518<=Vr;
XbG_H519<=Vr;
XbG_H52<=Vr;
XbG_H520<=Vr;
XbG_H521<=Vr;
XbG_H522<=Vr;
XbG_H523<=Vr;
XbG_H524<=Vr;
XbG_H525<=Vr;
XbG_H526<=Vr;
XbG_H527<=Vr;
XbG_H528<=Vr;
XbG_H529<=Vr;
XbG_H53<=Vr;
XbG_H530<=Vr;
XbG_H531<=Vr;
XbG_H532<=Vr;
XbG_H533<=Vr;
XbG_H534<=Vr;
XbG_H535<=Vr;
XbG_H536<=Vr;
XbG_H537<=Vr;
XbG_H538<=Vr;
XbG_H539<=Vr;
XbG_H54<=Vr;
XbG_H540<=Vr;
XbG_H541<=Vr;
XbG_H542<=Vr;
XbG_H543<=Vr;
XbG_H544<=Vr;
XbG_H545<=Vr;
XbG_H546<=Vr;
XbG_H547<=Vr;
XbG_H548<=Vr;
XbG_H549<=Vr;
XbG_H55<=Vr;
XbG_H550<=Vr;
XbG_H551<=Vr;
XbG_H552<=Vr;
XbG_H553<=Vr;
XbG_H554<=Vr;
XbG_H555<=Vr;
XbG_H556<=Vr;
XbG_H557<=Vr;
XbG_H558<=Vr;
XbG_H559<=Vr;
XbG_H56<=Vr;
XbG_H560<=Vr;
XbG_H561<=Vr;
XbG_H562<=Vr;
XbG_H563<=Vr;
XbG_H564<=Vr;
XbG_H565<=Vr;
XbG_H566<=Vr;
XbG_H567<=Vr;
XbG_H568<=Vr;
XbG_H569<=Vr;
XbG_H57<=Vr;
XbG_H570<=Vr;
XbG_H571<=Vr;
XbG_H572<=Vr;
XbG_H573<=Vr;
XbG_H574<=Vr;
XbG_H575<=Vr;
XbG_H576<=Vr;
XbG_H577<=Vr;
XbG_H578<=Vr;
XbG_H579<=Vr;
XbG_H58<=Vr;
XbG_H580<=Vr;
XbG_H581<=Vr;
XbG_H582<=Vr;
XbG_H583<=Vr;
XbG_H584<=Vr;
XbG_H585<=Vr;
XbG_H586<=Vr;
XbG_H587<=Vr;
XbG_H588<=Vr;
XbG_H589<=Vr;
XbG_H59<=Vr;
XbG_H590<=Vr;
XbG_H591<=Vr;
XbG_H592<=Vr;
XbG_H593<=Vr;
XbG_H594<=Vr;
XbG_H595<=Vr;
XbG_H596<=Vr;
XbG_H597<=Vr;
XbG_H598<=Vr;
XbG_H599<=Vr;
XbG_H6<=Vr;
XbG_H60<=Vr;
XbG_H600<=Vr;
XbG_H601<=Vr;
XbG_H602<=Vr;
XbG_H603<=Vr;
XbG_H604<=Vr;
XbG_H605<=Vr;
XbG_H606<=Vr;
XbG_H607<=Vr;
XbG_H608<=Vr;
XbG_H609<=Vr;
XbG_H61<=Vr;
XbG_H610<=Vr;
XbG_H611<=Vr;
XbG_H612<=Vr;
XbG_H613<=Vr;
XbG_H614<=Vr;
XbG_H615<=Vr;
XbG_H616<=Vr;
XbG_H617<=Vr;
XbG_H618<=Vr;
XbG_H619<=Vr;
XbG_H62<=Vr;
XbG_H620<=Vr;
XbG_H621<=Vr;
XbG_H622<=Vr;
XbG_H623<=Vr;
XbG_H624<=Vr;
XbG_H625<=Vr;
XbG_H626<=Vr;
XbG_H627<=Vr;
XbG_H628<=Vr;
XbG_H629<=Vr;
XbG_H63<=Vr;
XbG_H630<=Vr;
XbG_H631<=Vr;
XbG_H632<=Vr;
XbG_H633<=Vr;
XbG_H634<=Vr;
XbG_H635<=Vr;
XbG_H636<=Vr;
XbG_H637<=Vr;
XbG_H638<=Vr;
XbG_H639<=Vr;
XbG_H64<=Vr;
XbG_H640<=Vr;
XbG_H641<=Vr;
XbG_H642<=Vr;
XbG_H643<=Vr;
XbG_H644<=Vr;
XbG_H645<=Vr;
XbG_H646<=Vr;
XbG_H647<=Vr;
XbG_H648<=Vr;
XbG_H649<=Vr;
XbG_H65<=Vr;
XbG_H650<=Vr;
XbG_H651<=Vr;
XbG_H652<=Vr;
XbG_H653<=Vr;
XbG_H654<=Vr;
XbG_H655<=Vr;
XbG_H656<=Vr;
XbG_H657<=Vr;
XbG_H658<=Vr;
XbG_H659<=Vr;
XbG_H66<=Vr;
XbG_H660<=Vr;
XbG_H661<=(others=>'Z');
XbG_H662<=(others=>'Z');
XbG_H663<=(others=>'Z');
XbG_H664<=(others=>'Z');
XbG_H665<=(others=>'Z');
XbG_H666<=(others=>'Z');
XbG_H667<=(others=>'Z');
XbG_H668<=(others=>'Z');
XbG_H669<=(others=>'Z');
XbG_H67<=Vr;
XbG_H670<=(others=>'Z');
XbG_H671<=(others=>'Z');
XbG_H672<=(others=>'Z');
XbG_H673<=(others=>'Z');
XbG_H674<=(others=>'Z');
XbG_H675<=(others=>'Z');
XbG_H676<=(others=>'Z');
XbG_H677<=(others=>'Z');
XbG_H678<=(others=>'Z');
XbG_H679<=(others=>'Z');
XbG_H68<=Vr;
XbG_H680<=(others=>'Z');
XbG_H681<=(others=>'Z');
XbG_H682<=(others=>'Z');
XbG_H683<=(others=>'Z');
XbG_H684<=(others=>'Z');
XbG_H685<=(others=>'Z');
XbG_H686<=(others=>'Z');
XbG_H687<=(others=>'Z');
XbG_H688<=(others=>'Z');
XbG_H689<=(others=>'Z');
XbG_H69<=Vr;
XbG_H690<=(others=>'Z');
XbG_H691<=(others=>'Z');
XbG_H692<=(others=>'Z');
XbG_H693<=(others=>'Z');
XbG_H694<=(others=>'Z');
XbG_H695<=(others=>'Z');
XbG_H696<=(others=>'Z');
XbG_H697<=(others=>'Z');
XbG_H698<=(others=>'Z');
XbG_H699<=(others=>'Z');
XbG_H7<=Vr;
XbG_H70<=Vr;
XbG_H700<=(others=>'Z');
XbG_H701<=(others=>'Z');
XbG_H702<=(others=>'Z');
XbG_H703<=(others=>'Z');
XbG_H704<=(others=>'Z');
XbG_H705<=(others=>'Z');
XbG_H706<=(others=>'Z');
XbG_H707<=(others=>'Z');
XbG_H708<=(others=>'Z');
XbG_H709<=(others=>'Z');
XbG_H71<=Vr;
XbG_H710<=(others=>'Z');
XbG_H711<=(others=>'Z');
XbG_H712<=(others=>'Z');
XbG_H713<=(others=>'Z');
XbG_H714<=(others=>'Z');
XbG_H715<=(others=>'Z');
XbG_H716<=(others=>'Z');
XbG_H717<=(others=>'Z');
XbG_H718<=(others=>'Z');
XbG_H719<=(others=>'Z');
XbG_H72<=Vr;
XbG_H720<=(others=>'Z');
XbG_H721<=(others=>'Z');
XbG_H722<=Vr;
XbG_H723<=Vr;
XbG_H724<=Vr;
XbG_H725<=Vr;
XbG_H726<=Vr;
XbG_H727<=Vr;
XbG_H728<=Vr;
XbG_H729<=Vr;
XbG_H73<=Vr;
XbG_H730<=Vr;
XbG_H731<=Vr;
XbG_H732<=Vr;
XbG_H733<=Vr;
XbG_H734<=Vr;
XbG_H735<=Vr;
XbG_H74<=Vr;
XbG_H75<=Vr;
XbG_H76<=Vr;
XbG_H77<=Vr;
XbG_H78<=Vr;
XbG_H79<=Vr;
XbG_H8<=Vr;
XbG_H80<=Vr;
XbG_H81<=Vr;
XbG_H82<=Vr;
XbG_H83<=Vr;
XbG_H84<=Vr;
XbG_H85<=Vr;
XbG_H86<=Vr;
XbG_H87<=Vr;
XbG_H88<=Vr;
XbG_H89<=Vr;
XbG_H9<=Vr;
XbG_H90<=Vr;
XbG_H91<=Vr;
XbG_H92<=Vr;
XbG_H93<=Vr;
XbG_H94<=Vr;
XbG_H95<=Vr;
XbG_H96<=Vr;
XbG_H97<=Vr;
XbG_H98<=Vr;
XbG_H99<=Vr;
XbG_V0<=Vr;
XbG_V1<=Vr;
XbG_V10<=Vr;
XbG_V100<=Vw;
XbG_V101<=Vr;
XbG_V102<=Vw;
XbG_V103<=Vr;
XbG_V104<=Vw;
XbG_V105<=Vr;
XbG_V106<=Vw;
XbG_V107<=Vr;
XbG_V108<=Vw;
XbG_V109<=Vr;
XbG_V11<=Vr;
XbG_V110<=Vw;
XbG_V111<=Vr;
XbG_V112<=Vw;
XbG_V113<=Vr;
XbG_V114<=Vw;
XbG_V115<=Vr;
XbG_V116<=Vw;
XbG_V117<=Vr;
XbG_V118<=Vw;
XbG_V119<=Vr;
XbG_V12<=Vr;
XbG_V120<=Vw;
XbG_V121<=Vr;
XbG_V122<=Vw;
XbG_V123<=Vr;
XbG_V124<=Vw;
XbG_V125<=Vr;
XbG_V126<=Vw;
XbG_V127<=Vr;
XbG_V128<=Vw;
XbG_V129<=Vr;
XbG_V13<=Vr;
XbG_V130<=Vw;
XbG_V131<=Vr;
XbG_V132<=Vw;
XbG_V133<=Vr;
XbG_V134<=Vw;
XbG_V135<=Vr;
XbG_V136<=Vw;
XbG_V137<=Vr;
XbG_V138<=Vw;
XbG_V139<=Vr;
XbG_V14<=Vr;
XbG_V140<=Vw;
XbG_V141<=Vr;
XbG_V142<=Vw;
XbG_V143<=Vr;
XbG_V144<=Vw;
XbG_V145<=Vr;
XbG_V146<=Vw;
XbG_V147<=Vr;
XbG_V148<=Vw;
XbG_V149<=Vr;
XbG_V15<=Vr;
XbG_V150<=Vw;
XbG_V151<=Vr;
XbG_V152<=Vw;
XbG_V153<=Vr;
XbG_V154<=Vw;
XbG_V155<=Vr;
XbG_V156<=Vw;
XbG_V157<=Vr;
XbG_V158<=Vw;
XbG_V159<=Vr;
XbG_V16<=Vr;
XbG_V160<=Vw;
XbG_V161<=Vr;
XbG_V162<=Vw;
XbG_V163<=Vr;
XbG_V164<=Vw;
XbG_V165<=Vr;
XbG_V166<=Vw;
XbG_V167<=Vr;
XbG_V168<=Vw;
XbG_V169<=Vr;
XbG_V17<=Vr;
XbG_V170<=Vw;
XbG_V171<=Vr;
XbG_V172<=Vw;
XbG_V173<=Vr;
XbG_V174<=Vw;
XbG_V175<=Vr;
XbG_V176<=Vw;
XbG_V177<=Vr;
XbG_V178<=Vw;
XbG_V179<=Vr;
XbG_V18<=Vr;
XbG_V180<=Vw;
XbG_V181<=Vr;
XbG_V182<=Vw;
XbG_V183<=Vr;
XbG_V184<=Vw;
XbG_V185<=Vr;
XbG_V186<=Vw;
XbG_V187<=Vr;
XbG_V188<=Vw;
XbG_V189<=Vr;
XbG_V19<=Vr;
XbG_V2<=Vr;
XbG_V20<=Vr;
XbG_V21<=Vr;
XbG_V22<=Vr;
XbG_V23<=Vr;
XbG_V24<=Vr;
XbG_V25<=Vr;
XbG_V26<=Vr;
XbG_V27<=Vr;
XbG_V28<=Vr;
XbG_V29<=Vr;
XbG_V3<=Vr;
XbG_V30<=Vr;
XbG_V31<=Vr;
XbG_V32<=Vr;
XbG_V33<=Vr;
XbG_V34<=Vr;
XbG_V35<=Vr;
XbG_V36<=Vr;
XbG_V37<=Vr;
XbG_V38<=Vr;
XbG_V39<=Vr;
XbG_V4<=Vr;
XbG_V40<=Vr;
XbG_V41<=Vr;
XbG_V42<=Vr;
XbG_V43<=Vr;
XbG_V44<=Vr;
XbG_V45<=Vr;
XbG_V46<=Vr;
XbG_V47<=Vr;
XbG_V48<=Vr;
XbG_V49<=Vr;
XbG_V5<=Vr;
XbG_V50<=Vr;
XbG_V51<=Vr;
XbG_V52<=Vr;
XbG_V53<=Vr;
XbG_V54<=Vr;
XbG_V55<=Vr;
XbG_V56<=Vr;
XbG_V57<=Vr;
XbG_V58<=Vr;
XbG_V59<=Vr;
XbG_V6<=Vr;
XbG_V60<=Vr;
XbG_V61<=Vr;
XbG_V62<=Vr;
XbG_V63<=Vr;
XbG_V64<=Vr;
XbG_V65<=Vr;
XbG_V66<=Vr;
XbG_V67<=Vr;
XbG_V68<=Vw;
XbG_V69<=Vr;
XbG_V7<=Vr;
XbG_V70<=Vw;
XbG_V71<=Vr;
XbG_V72<=Vw;
XbG_V73<=Vr;
XbG_V74<=Vw;
XbG_V75<=Vr;
XbG_V76<=Vw;
XbG_V77<=Vr;
XbG_V78<=Vw;
XbG_V79<=Vr;
XbG_V8<=Vr;
XbG_V80<=Vw;
XbG_V81<=Vr;
XbG_V82<=Vw;
XbG_V83<=Vr;
XbG_V84<=Vw;
XbG_V85<=Vr;
XbG_V86<=Vw;
XbG_V87<=Vr;
XbG_V88<=Vw;
XbG_V89<=Vr;
XbG_V9<=Vr;
XbG_V90<=Vw;
XbG_V91<=Vr;
XbG_V92<=Vw;
XbG_V93<=Vr;
XbG_V94<=Vw;
XbG_V95<=Vr;
XbG_V96<=Vw;
XbG_V97<=Vr;
XbG_V98<=Vw;
XbG_V99<=Vr;

next_state<=G_SS;

when G_SS =>

XbG_H0<=Vr;
XbG_H1<=(others=>'Z');
XbG_H10<=(others=>'Z');
XbG_H100<=(others=>'Z');
XbG_H101<=(others=>'Z');
XbG_H102<=(others=>'Z');
XbG_H103<=(others=>'Z');
XbG_H104<=(others=>'Z');
XbG_H105<=(others=>'Z');
XbG_H106<=(others=>'Z');
XbG_H107<=(others=>'Z');
XbG_H108<=(others=>'Z');
XbG_H109<=(others=>'Z');
XbG_H11<=(others=>'Z');
XbG_H110<=(others=>'Z');
XbG_H111<=(others=>'Z');
XbG_H112<=(others=>'Z');
XbG_H113<=(others=>'Z');
XbG_H114<=(others=>'Z');
XbG_H115<=(others=>'Z');
XbG_H116<=(others=>'Z');
XbG_H117<=(others=>'Z');
XbG_H118<=(others=>'Z');
XbG_H119<=(others=>'Z');
XbG_H12<=(others=>'Z');
XbG_H120<=(others=>'Z');
XbG_H121<=(others=>'Z');
XbG_H122<=(others=>'Z');
XbG_H123<=(others=>'Z');
XbG_H124<=(others=>'Z');
XbG_H125<=(others=>'Z');
XbG_H126<=(others=>'Z');
XbG_H127<=(others=>'Z');
XbG_H128<=(others=>'Z');
XbG_H129<=(others=>'Z');
XbG_H13<=(others=>'Z');
XbG_H130<=(others=>'Z');
XbG_H131<=(others=>'Z');
XbG_H132<=(others=>'Z');
XbG_H133<=(others=>'Z');
XbG_H134<=(others=>'Z');
XbG_H135<=(others=>'Z');
XbG_H136<=(others=>'Z');
XbG_H137<=(others=>'Z');
XbG_H138<=(others=>'Z');
XbG_H139<=(others=>'Z');
XbG_H14<=(others=>'Z');
XbG_H140<=(others=>'Z');
XbG_H141<=(others=>'Z');
XbG_H142<=(others=>'Z');
XbG_H143<=(others=>'Z');
XbG_H144<=(others=>'Z');
XbG_H145<=(others=>'Z');
XbG_H146<=(others=>'Z');
XbG_H147<=(others=>'Z');
XbG_H148<=(others=>'Z');
XbG_H149<=(others=>'Z');
XbG_H15<=(others=>'Z');
XbG_H150<=(others=>'Z');
XbG_H151<=(others=>'Z');
XbG_H152<=(others=>'Z');
XbG_H153<=(others=>'Z');
XbG_H154<=(others=>'Z');
XbG_H155<=(others=>'Z');
XbG_H156<=(others=>'Z');
XbG_H157<=(others=>'Z');
XbG_H158<=(others=>'Z');
XbG_H159<=(others=>'Z');
XbG_H16<=(others=>'Z');
XbG_H160<=(others=>'Z');
XbG_H161<=(others=>'Z');
XbG_H162<=(others=>'Z');
XbG_H163<=(others=>'Z');
XbG_H164<=(others=>'Z');
XbG_H165<=(others=>'Z');
XbG_H166<=(others=>'Z');
XbG_H167<=(others=>'Z');
XbG_H168<=(others=>'Z');
XbG_H169<=(others=>'Z');
XbG_H17<=(others=>'Z');
XbG_H170<=(others=>'Z');
XbG_H171<=(others=>'Z');
XbG_H172<=(others=>'Z');
XbG_H173<=(others=>'Z');
XbG_H174<=(others=>'Z');
XbG_H175<=(others=>'Z');
XbG_H176<=(others=>'Z');
XbG_H177<=(others=>'Z');
XbG_H178<=(others=>'Z');
XbG_H179<=(others=>'Z');
XbG_H18<=(others=>'Z');
XbG_H180<=(others=>'Z');
XbG_H181<=(others=>'Z');
XbG_H182<=(others=>'Z');
XbG_H183<=(others=>'Z');
XbG_H184<=(others=>'Z');
XbG_H185<=(others=>'Z');
XbG_H186<=(others=>'Z');
XbG_H187<=(others=>'Z');
XbG_H188<=(others=>'Z');
XbG_H189<=(others=>'Z');
XbG_H19<=(others=>'Z');
XbG_H190<=(others=>'Z');
XbG_H191<=(others=>'Z');
XbG_H192<=(others=>'Z');
XbG_H193<=(others=>'Z');
XbG_H194<=(others=>'Z');
XbG_H195<=(others=>'Z');
XbG_H196<=(others=>'Z');
XbG_H197<=(others=>'Z');
XbG_H198<=(others=>'Z');
XbG_H199<=(others=>'Z');
XbG_H2<=(others=>'Z');
XbG_H20<=(others=>'Z');
XbG_H200<=(others=>'Z');
XbG_H201<=(others=>'Z');
XbG_H202<=(others=>'Z');
XbG_H203<=(others=>'Z');
XbG_H204<=(others=>'Z');
XbG_H205<=(others=>'Z');
XbG_H206<=(others=>'Z');
XbG_H207<=(others=>'Z');
XbG_H208<=(others=>'Z');
XbG_H209<=(others=>'Z');
XbG_H21<=(others=>'Z');
XbG_H210<=(others=>'Z');
XbG_H211<=(others=>'Z');
XbG_H212<=(others=>'Z');
XbG_H213<=(others=>'Z');
XbG_H214<=(others=>'Z');
XbG_H215<=(others=>'Z');
XbG_H216<=(others=>'Z');
XbG_H217<=(others=>'Z');
XbG_H218<=(others=>'Z');
XbG_H219<=(others=>'Z');
XbG_H22<=(others=>'Z');
XbG_H220<=(others=>'Z');
XbG_H221<=(others=>'Z');
XbG_H222<=(others=>'Z');
XbG_H223<=(others=>'Z');
XbG_H224<=(others=>'Z');
XbG_H225<=(others=>'Z');
XbG_H226<=(others=>'Z');
XbG_H227<=(others=>'Z');
XbG_H228<=(others=>'Z');
XbG_H229<=(others=>'Z');
XbG_H23<=(others=>'Z');
XbG_H230<=(others=>'Z');
XbG_H231<=(others=>'Z');
XbG_H232<=(others=>'Z');
XbG_H233<=(others=>'Z');
XbG_H234<=(others=>'Z');
XbG_H235<=(others=>'Z');
XbG_H236<=(others=>'Z');
XbG_H237<=(others=>'Z');
XbG_H238<=(others=>'Z');
XbG_H239<=(others=>'Z');
XbG_H24<=(others=>'Z');
XbG_H240<=(others=>'Z');
XbG_H241<=(others=>'Z');
XbG_H242<=(others=>'Z');
XbG_H243<=(others=>'Z');
XbG_H244<=(others=>'Z');
XbG_H245<=(others=>'Z');
XbG_H246<=(others=>'Z');
XbG_H247<=(others=>'Z');
XbG_H248<=(others=>'Z');
XbG_H249<=(others=>'Z');
XbG_H25<=(others=>'Z');
XbG_H250<=(others=>'Z');
XbG_H251<=(others=>'Z');
XbG_H252<=(others=>'Z');
XbG_H253<=(others=>'Z');
XbG_H254<=(others=>'Z');
XbG_H255<=(others=>'Z');
XbG_H256<=(others=>'Z');
XbG_H257<=(others=>'Z');
XbG_H258<=(others=>'Z');
XbG_H259<=(others=>'Z');
XbG_H26<=(others=>'Z');
XbG_H260<=(others=>'Z');
XbG_H261<=(others=>'Z');
XbG_H262<=(others=>'Z');
XbG_H263<=(others=>'Z');
XbG_H264<=(others=>'Z');
XbG_H265<=(others=>'Z');
XbG_H266<=(others=>'Z');
XbG_H267<=(others=>'Z');
XbG_H268<=(others=>'Z');
XbG_H269<=(others=>'Z');
XbG_H27<=(others=>'Z');
XbG_H270<=(others=>'Z');
XbG_H271<=(others=>'Z');
XbG_H272<=(others=>'Z');
XbG_H273<=(others=>'Z');
XbG_H274<=(others=>'Z');
XbG_H275<=(others=>'Z');
XbG_H276<=(others=>'Z');
XbG_H277<=(others=>'Z');
XbG_H278<=(others=>'Z');
XbG_H279<=(others=>'Z');
XbG_H28<=(others=>'Z');
XbG_H280<=(others=>'Z');
XbG_H281<=(others=>'Z');
XbG_H282<=(others=>'Z');
XbG_H283<=(others=>'Z');
XbG_H284<=(others=>'Z');
XbG_H285<=(others=>'Z');
XbG_H286<=(others=>'Z');
XbG_H287<=(others=>'Z');
XbG_H288<=(others=>'Z');
XbG_H289<=(others=>'Z');
XbG_H29<=(others=>'Z');
XbG_H290<=(others=>'Z');
XbG_H291<=(others=>'Z');
XbG_H292<=(others=>'Z');
XbG_H293<=(others=>'Z');
XbG_H294<=(others=>'Z');
XbG_H295<=(others=>'Z');
XbG_H296<=(others=>'Z');
XbG_H297<=(others=>'Z');
XbG_H298<=(others=>'Z');
XbG_H299<=(others=>'Z');
XbG_H3<=(others=>'Z');
XbG_H30<=(others=>'Z');
XbG_H300<=(others=>'Z');
XbG_H301<=(others=>'Z');
XbG_H302<=(others=>'Z');
XbG_H303<=(others=>'Z');
XbG_H304<=(others=>'Z');
XbG_H305<=(others=>'Z');
XbG_H306<=(others=>'Z');
XbG_H307<=(others=>'Z');
XbG_H308<=(others=>'Z');
XbG_H309<=(others=>'Z');
XbG_H31<=(others=>'Z');
XbG_H310<=(others=>'Z');
XbG_H311<=(others=>'Z');
XbG_H312<=(others=>'Z');
XbG_H313<=(others=>'Z');
XbG_H314<=(others=>'Z');
XbG_H315<=(others=>'Z');
XbG_H316<=(others=>'Z');
XbG_H317<=(others=>'Z');
XbG_H318<=(others=>'Z');
XbG_H319<=(others=>'Z');
XbG_H32<=(others=>'Z');
XbG_H320<=(others=>'Z');
XbG_H321<=(others=>'Z');
XbG_H322<=(others=>'Z');
XbG_H323<=(others=>'Z');
XbG_H324<=(others=>'Z');
XbG_H325<=(others=>'Z');
XbG_H326<=(others=>'Z');
XbG_H327<=(others=>'Z');
XbG_H328<=(others=>'Z');
XbG_H329<=(others=>'Z');
XbG_H33<=(others=>'Z');
XbG_H330<=(others=>'Z');
XbG_H331<=(others=>'Z');
XbG_H332<=(others=>'Z');
XbG_H333<=(others=>'Z');
XbG_H334<=(others=>'Z');
XbG_H335<=(others=>'Z');
XbG_H336<=(others=>'Z');
XbG_H337<=(others=>'Z');
XbG_H338<=(others=>'Z');
XbG_H339<=(others=>'Z');
XbG_H34<=(others=>'Z');
XbG_H340<=(others=>'Z');
XbG_H341<=(others=>'Z');
XbG_H342<=(others=>'Z');
XbG_H343<=(others=>'Z');
XbG_H344<=(others=>'Z');
XbG_H345<=(others=>'Z');
XbG_H346<=(others=>'Z');
XbG_H347<=(others=>'Z');
XbG_H348<=(others=>'Z');
XbG_H349<=(others=>'Z');
XbG_H35<=(others=>'Z');
XbG_H350<=(others=>'Z');
XbG_H351<=(others=>'Z');
XbG_H352<=(others=>'Z');
XbG_H353<=(others=>'Z');
XbG_H354<=(others=>'Z');
XbG_H355<=(others=>'Z');
XbG_H356<=(others=>'Z');
XbG_H357<=(others=>'Z');
XbG_H358<=(others=>'Z');
XbG_H359<=(others=>'Z');
XbG_H36<=(others=>'Z');
XbG_H360<=(others=>'Z');
XbG_H361<=(others=>'Z');
XbG_H362<=(others=>'Z');
XbG_H363<=(others=>'Z');
XbG_H364<=(others=>'Z');
XbG_H365<=(others=>'Z');
XbG_H366<=(others=>'Z');
XbG_H367<=(others=>'Z');
XbG_H368<=(others=>'Z');
XbG_H369<=(others=>'Z');
XbG_H37<=(others=>'Z');
XbG_H370<=(others=>'Z');
XbG_H371<=(others=>'Z');
XbG_H372<=(others=>'Z');
XbG_H373<=(others=>'Z');
XbG_H374<=(others=>'Z');
XbG_H375<=(others=>'Z');
XbG_H376<=(others=>'Z');
XbG_H377<=(others=>'Z');
XbG_H378<=(others=>'Z');
XbG_H379<=(others=>'Z');
XbG_H38<=(others=>'Z');
XbG_H380<=(others=>'Z');
XbG_H381<=(others=>'Z');
XbG_H382<=(others=>'Z');
XbG_H383<=(others=>'Z');
XbG_H384<=(others=>'Z');
XbG_H385<=(others=>'Z');
XbG_H386<=(others=>'Z');
XbG_H387<=(others=>'Z');
XbG_H388<=(others=>'Z');
XbG_H389<=(others=>'Z');
XbG_H39<=(others=>'Z');
XbG_H390<=(others=>'Z');
XbG_H391<=(others=>'Z');
XbG_H392<=(others=>'Z');
XbG_H393<=(others=>'Z');
XbG_H394<=(others=>'Z');
XbG_H395<=(others=>'Z');
XbG_H396<=(others=>'Z');
XbG_H397<=(others=>'Z');
XbG_H398<=(others=>'Z');
XbG_H399<=(others=>'Z');
XbG_H4<=(others=>'Z');
XbG_H40<=(others=>'Z');
XbG_H400<=(others=>'Z');
XbG_H401<=(others=>'Z');
XbG_H402<=(others=>'Z');
XbG_H403<=(others=>'Z');
XbG_H404<=(others=>'Z');
XbG_H405<=(others=>'Z');
XbG_H406<=(others=>'Z');
XbG_H407<=(others=>'Z');
XbG_H408<=(others=>'Z');
XbG_H409<=(others=>'Z');
XbG_H41<=(others=>'Z');
XbG_H410<=(others=>'Z');
XbG_H411<=(others=>'Z');
XbG_H412<=(others=>'Z');
XbG_H413<=(others=>'Z');
XbG_H414<=(others=>'Z');
XbG_H415<=(others=>'Z');
XbG_H416<=(others=>'Z');
XbG_H417<=(others=>'Z');
XbG_H418<=(others=>'Z');
XbG_H419<=(others=>'Z');
XbG_H42<=(others=>'Z');
XbG_H420<=(others=>'Z');
XbG_H421<=(others=>'Z');
XbG_H422<=(others=>'Z');
XbG_H423<=(others=>'Z');
XbG_H424<=(others=>'Z');
XbG_H425<=(others=>'Z');
XbG_H426<=(others=>'Z');
XbG_H427<=(others=>'Z');
XbG_H428<=(others=>'Z');
XbG_H429<=(others=>'Z');
XbG_H43<=(others=>'Z');
XbG_H430<=(others=>'Z');
XbG_H431<=(others=>'Z');
XbG_H432<=(others=>'Z');
XbG_H433<=(others=>'Z');
XbG_H434<=(others=>'Z');
XbG_H435<=(others=>'Z');
XbG_H436<=(others=>'Z');
XbG_H437<=(others=>'Z');
XbG_H438<=(others=>'Z');
XbG_H439<=(others=>'Z');
XbG_H44<=(others=>'Z');
XbG_H440<=(others=>'Z');
XbG_H441<=(others=>'Z');
XbG_H442<=(others=>'Z');
XbG_H443<=(others=>'Z');
XbG_H444<=(others=>'Z');
XbG_H445<=(others=>'Z');
XbG_H446<=(others=>'Z');
XbG_H447<=(others=>'Z');
XbG_H448<=(others=>'Z');
XbG_H449<=(others=>'Z');
XbG_H45<=(others=>'Z');
XbG_H450<=(others=>'Z');
XbG_H451<=(others=>'Z');
XbG_H452<=(others=>'Z');
XbG_H453<=(others=>'Z');
XbG_H454<=(others=>'Z');
XbG_H455<=(others=>'Z');
XbG_H456<=(others=>'Z');
XbG_H457<=(others=>'Z');
XbG_H458<=(others=>'Z');
XbG_H459<=(others=>'Z');
XbG_H46<=(others=>'Z');
XbG_H460<=(others=>'Z');
XbG_H461<=(others=>'Z');
XbG_H462<=(others=>'Z');
XbG_H463<=(others=>'Z');
XbG_H464<=(others=>'Z');
XbG_H465<=(others=>'Z');
XbG_H466<=(others=>'Z');
XbG_H467<=(others=>'Z');
XbG_H468<=(others=>'Z');
XbG_H469<=(others=>'Z');
XbG_H47<=(others=>'Z');
XbG_H470<=(others=>'Z');
XbG_H471<=(others=>'Z');
XbG_H472<=(others=>'Z');
XbG_H473<=(others=>'Z');
XbG_H474<=(others=>'Z');
XbG_H475<=(others=>'Z');
XbG_H476<=(others=>'Z');
XbG_H477<=(others=>'Z');
XbG_H478<=(others=>'Z');
XbG_H479<=(others=>'Z');
XbG_H48<=(others=>'Z');
XbG_H480<=(others=>'Z');
XbG_H481<=(others=>'Z');
XbG_H482<=(others=>'Z');
XbG_H483<=(others=>'Z');
XbG_H484<=(others=>'Z');
XbG_H485<=(others=>'Z');
XbG_H486<=(others=>'Z');
XbG_H487<=(others=>'Z');
XbG_H488<=(others=>'Z');
XbG_H489<=(others=>'Z');
XbG_H49<=(others=>'Z');
XbG_H490<=(others=>'Z');
XbG_H491<=(others=>'Z');
XbG_H492<=(others=>'Z');
XbG_H493<=(others=>'Z');
XbG_H494<=(others=>'Z');
XbG_H495<=(others=>'Z');
XbG_H496<=(others=>'Z');
XbG_H497<=(others=>'Z');
XbG_H498<=(others=>'Z');
XbG_H499<=(others=>'Z');
XbG_H5<=(others=>'Z');
XbG_H50<=(others=>'Z');
XbG_H500<=(others=>'Z');
XbG_H501<=(others=>'Z');
XbG_H502<=(others=>'Z');
XbG_H503<=(others=>'Z');
XbG_H504<=(others=>'Z');
XbG_H505<=(others=>'Z');
XbG_H506<=(others=>'Z');
XbG_H507<=(others=>'Z');
XbG_H508<=(others=>'Z');
XbG_H509<=(others=>'Z');
XbG_H51<=(others=>'Z');
XbG_H510<=(others=>'Z');
XbG_H511<=(others=>'Z');
XbG_H512<=(others=>'Z');
XbG_H513<=(others=>'Z');
XbG_H514<=(others=>'Z');
XbG_H515<=(others=>'Z');
XbG_H516<=(others=>'Z');
XbG_H517<=(others=>'Z');
XbG_H518<=(others=>'Z');
XbG_H519<=(others=>'Z');
XbG_H52<=(others=>'Z');
XbG_H520<=(others=>'Z');
XbG_H521<=(others=>'Z');
XbG_H522<=(others=>'Z');
XbG_H523<=(others=>'Z');
XbG_H524<=(others=>'Z');
XbG_H525<=(others=>'Z');
XbG_H526<=(others=>'Z');
XbG_H527<=(others=>'Z');
XbG_H528<=(others=>'Z');
XbG_H529<=(others=>'Z');
XbG_H53<=(others=>'Z');
XbG_H530<=(others=>'Z');
XbG_H531<=(others=>'Z');
XbG_H532<=(others=>'Z');
XbG_H533<=(others=>'Z');
XbG_H534<=(others=>'Z');
XbG_H535<=(others=>'Z');
XbG_H536<=(others=>'Z');
XbG_H537<=(others=>'Z');
XbG_H538<=(others=>'Z');
XbG_H539<=(others=>'Z');
XbG_H54<=(others=>'Z');
XbG_H540<=(others=>'Z');
XbG_H541<=(others=>'Z');
XbG_H542<=(others=>'Z');
XbG_H543<=(others=>'Z');
XbG_H544<=(others=>'Z');
XbG_H545<=(others=>'Z');
XbG_H546<=(others=>'Z');
XbG_H547<=(others=>'Z');
XbG_H548<=(others=>'Z');
XbG_H549<=(others=>'Z');
XbG_H55<=(others=>'Z');
XbG_H550<=(others=>'Z');
XbG_H551<=(others=>'Z');
XbG_H552<=(others=>'Z');
XbG_H553<=(others=>'Z');
XbG_H554<=(others=>'Z');
XbG_H555<=(others=>'Z');
XbG_H556<=(others=>'Z');
XbG_H557<=(others=>'Z');
XbG_H558<=(others=>'Z');
XbG_H559<=(others=>'Z');
XbG_H56<=(others=>'Z');
XbG_H560<=(others=>'Z');
XbG_H561<=(others=>'Z');
XbG_H562<=(others=>'Z');
XbG_H563<=(others=>'Z');
XbG_H564<=(others=>'Z');
XbG_H565<=(others=>'Z');
XbG_H566<=(others=>'Z');
XbG_H567<=(others=>'Z');
XbG_H568<=(others=>'Z');
XbG_H569<=(others=>'Z');
XbG_H57<=(others=>'Z');
XbG_H570<=(others=>'Z');
XbG_H571<=(others=>'Z');
XbG_H572<=(others=>'Z');
XbG_H573<=(others=>'Z');
XbG_H574<=(others=>'Z');
XbG_H575<=(others=>'Z');
XbG_H576<=(others=>'Z');
XbG_H577<=(others=>'Z');
XbG_H578<=(others=>'Z');
XbG_H579<=(others=>'Z');
XbG_H58<=(others=>'Z');
XbG_H580<=(others=>'Z');
XbG_H581<=(others=>'Z');
XbG_H582<=(others=>'Z');
XbG_H583<=(others=>'Z');
XbG_H584<=(others=>'Z');
XbG_H585<=(others=>'Z');
XbG_H586<=(others=>'Z');
XbG_H587<=(others=>'Z');
XbG_H588<=(others=>'Z');
XbG_H589<=(others=>'Z');
XbG_H59<=(others=>'Z');
XbG_H590<=(others=>'Z');
XbG_H591<=(others=>'Z');
XbG_H592<=(others=>'Z');
XbG_H593<=(others=>'Z');
XbG_H594<=(others=>'Z');
XbG_H595<=(others=>'Z');
XbG_H596<=(others=>'Z');
XbG_H597<=(others=>'Z');
XbG_H598<=(others=>'Z');
XbG_H599<=(others=>'Z');
XbG_H6<=(others=>'Z');
XbG_H60<=(others=>'Z');
XbG_H600<=(others=>'Z');
XbG_H601<=(others=>'Z');
XbG_H602<=(others=>'Z');
XbG_H603<=(others=>'Z');
XbG_H604<=(others=>'Z');
XbG_H605<=(others=>'Z');
XbG_H606<=(others=>'Z');
XbG_H607<=(others=>'Z');
XbG_H608<=(others=>'Z');
XbG_H609<=(others=>'Z');
XbG_H61<=(others=>'Z');
XbG_H610<=(others=>'Z');
XbG_H611<=(others=>'Z');
XbG_H612<=(others=>'Z');
XbG_H613<=(others=>'Z');
XbG_H614<=(others=>'Z');
XbG_H615<=(others=>'Z');
XbG_H616<=(others=>'Z');
XbG_H617<=(others=>'Z');
XbG_H618<=(others=>'Z');
XbG_H619<=(others=>'Z');
XbG_H62<=(others=>'Z');
XbG_H620<=(others=>'Z');
XbG_H621<=(others=>'Z');
XbG_H622<=(others=>'Z');
XbG_H623<=(others=>'Z');
XbG_H624<=(others=>'Z');
XbG_H625<=(others=>'Z');
XbG_H626<=(others=>'Z');
XbG_H627<=(others=>'Z');
XbG_H628<=(others=>'Z');
XbG_H629<=(others=>'Z');
XbG_H63<=(others=>'Z');
XbG_H630<=(others=>'Z');
XbG_H631<=(others=>'Z');
XbG_H632<=(others=>'Z');
XbG_H633<=(others=>'Z');
XbG_H634<=(others=>'Z');
XbG_H635<=(others=>'Z');
XbG_H636<=(others=>'Z');
XbG_H637<=(others=>'Z');
XbG_H638<=(others=>'Z');
XbG_H639<=(others=>'Z');
XbG_H64<=(others=>'Z');
XbG_H640<=(others=>'Z');
XbG_H641<=(others=>'Z');
XbG_H642<=(others=>'Z');
XbG_H643<=(others=>'Z');
XbG_H644<=(others=>'Z');
XbG_H645<=(others=>'Z');
XbG_H646<=(others=>'Z');
XbG_H647<=(others=>'Z');
XbG_H648<=(others=>'Z');
XbG_H649<=(others=>'Z');
XbG_H65<=(others=>'Z');
XbG_H650<=(others=>'Z');
XbG_H651<=(others=>'Z');
XbG_H652<=(others=>'Z');
XbG_H653<=(others=>'Z');
XbG_H654<=(others=>'Z');
XbG_H655<=(others=>'Z');
XbG_H656<=(others=>'Z');
XbG_H657<=(others=>'Z');
XbG_H658<=(others=>'Z');
XbG_H659<=(others=>'Z');
XbG_H66<=(others=>'Z');
XbG_H660<=(others=>'Z');
XbG_H661<=Vw;
XbG_H662<=Vw;
XbG_H663<=Vw;
XbG_H664<=Vw;
XbG_H665<=Vw;
XbG_H666<=Vw;
XbG_H667<=Vw;
XbG_H668<=Vw;
XbG_H669<=Vw;
XbG_H67<=(others=>'Z');
XbG_H670<=Vw;
XbG_H671<=Vw;
XbG_H672<=Vw;
XbG_H673<=Vw;
XbG_H674<=Vw;
XbG_H675<=Vw;
XbG_H676<=Vw;
XbG_H677<=Vw;
XbG_H678<=Vw;
XbG_H679<=Vw;
XbG_H68<=(others=>'Z');
XbG_H680<=Vw;
XbG_H681<=Vw;
XbG_H682<=Vw;
XbG_H683<=Vw;
XbG_H684<=Vw;
XbG_H685<=Vw;
XbG_H686<=Vw;
XbG_H687<=Vw;
XbG_H688<=Vw;
XbG_H689<=Vw;
XbG_H69<=(others=>'Z');
XbG_H690<=Vw;
XbG_H691<=Vw;
XbG_H692<=Vw;
XbG_H693<=Vw;
XbG_H694<=Vw;
XbG_H695<=Vw;
XbG_H696<=Vw;
XbG_H697<=Vw;
XbG_H698<=Vw;
XbG_H699<=Vw;
XbG_H7<=(others=>'Z');
XbG_H70<=(others=>'Z');
XbG_H700<=Vw;
XbG_H701<=Vw;
XbG_H702<=Vw;
XbG_H703<=Vw;
XbG_H704<=Vw;
XbG_H705<=Vw;
XbG_H706<=Vw;
XbG_H707<=Vw;
XbG_H708<=Vw;
XbG_H709<=Vw;
XbG_H71<=(others=>'Z');
XbG_H710<=Vw;
XbG_H711<=Vw;
XbG_H712<=Vw;
XbG_H713<=Vw;
XbG_H714<=Vw;
XbG_H715<=Vw;
XbG_H716<=Vw;
XbG_H717<=Vw;
XbG_H718<=Vw;
XbG_H719<=Vw;
XbG_H72<=(others=>'Z');
XbG_H720<=Vw;
XbG_H721<=Vw;
XbG_H722<=zero;
XbG_H723<=zero;
XbG_H724<=zero;
XbG_H725<=zero;
XbG_H726<=zero;
XbG_H727<=zero;
XbG_H728<=zero;
XbG_H729<=zero;
XbG_H73<=(others=>'Z');
XbG_H730<=zero;
XbG_H731<=zero;
XbG_H732<=zero;
XbG_H733<=zero;
XbG_H734<=zero;
XbG_H735<=zero;
XbG_H74<=(others=>'Z');
XbG_H75<=(others=>'Z');
XbG_H76<=(others=>'Z');
XbG_H77<=(others=>'Z');
XbG_H78<=(others=>'Z');
XbG_H79<=(others=>'Z');
XbG_H8<=(others=>'Z');
XbG_H80<=(others=>'Z');
XbG_H81<=(others=>'Z');
XbG_H82<=(others=>'Z');
XbG_H83<=(others=>'Z');
XbG_H84<=(others=>'Z');
XbG_H85<=(others=>'Z');
XbG_H86<=(others=>'Z');
XbG_H87<=(others=>'Z');
XbG_H88<=(others=>'Z');
XbG_H89<=(others=>'Z');
XbG_H9<=(others=>'Z');
XbG_H90<=(others=>'Z');
XbG_H91<=(others=>'Z');
XbG_H92<=(others=>'Z');
XbG_H93<=(others=>'Z');
XbG_H94<=(others=>'Z');
XbG_H95<=(others=>'Z');
XbG_H96<=(others=>'Z');
XbG_H97<=(others=>'Z');
XbG_H98<=(others=>'Z');
XbG_H99<=(others=>'Z');
XbG_V0<=(others=>'Z');
XbG_V1<=(others=>'Z');
XbG_V10<=(others=>'Z');
XbG_V100<=Vr, (others=>'Z') after 1 ps;
XbG_V101<=(others=>'Z');
XbG_V102<=Vr, (others=>'Z') after 1 ps;
XbG_V103<=(others=>'Z');
XbG_V104<=Vr, (others=>'Z') after 1 ps;
XbG_V105<=(others=>'Z');
XbG_V106<=Vr, (others=>'Z') after 1 ps;
XbG_V107<=(others=>'Z');
XbG_V108<=Vr, (others=>'Z') after 1 ps;
XbG_V109<=(others=>'Z');
XbG_V11<=(others=>'Z');
XbG_V110<=Vr, (others=>'Z') after 1 ps;
XbG_V111<=(others=>'Z');
XbG_V112<=Vr, (others=>'Z') after 1 ps;
XbG_V113<=(others=>'Z');
XbG_V114<=Vr, (others=>'Z') after 1 ps;
XbG_V115<=(others=>'Z');
XbG_V116<=Vr, (others=>'Z') after 1 ps;
XbG_V117<=(others=>'Z');
XbG_V118<=Vr, (others=>'Z') after 1 ps;
XbG_V119<=(others=>'Z');
XbG_V12<=(others=>'Z');
XbG_V120<=Vr, (others=>'Z') after 1 ps;
XbG_V121<=(others=>'Z');
XbG_V122<=Vr, (others=>'Z') after 1 ps;
XbG_V123<=(others=>'Z');
XbG_V124<=Vr, (others=>'Z') after 1 ps;
XbG_V125<=(others=>'Z');
XbG_V126<=Vr, (others=>'Z') after 1 ps;
XbG_V127<=(others=>'Z');
XbG_V128<=Vr, (others=>'Z') after 1 ps;
XbG_V129<=(others=>'Z');
XbG_V13<=(others=>'Z');
XbG_V130<=Vr, (others=>'Z') after 1 ps;
XbG_V131<=(others=>'Z');
XbG_V132<=Vr, (others=>'Z') after 1 ps;
XbG_V133<=(others=>'Z');
XbG_V134<=Vr, (others=>'Z') after 1 ps;
XbG_V135<=(others=>'Z');
XbG_V136<=Vr, (others=>'Z') after 1 ps;
XbG_V137<=(others=>'Z');
XbG_V138<=Vr, (others=>'Z') after 1 ps;
XbG_V139<=(others=>'Z');
XbG_V14<=(others=>'Z');
XbG_V140<=Vr, (others=>'Z') after 1 ps;
XbG_V141<=(others=>'Z');
XbG_V142<=Vr, (others=>'Z') after 1 ps;
XbG_V143<=(others=>'Z');
XbG_V144<=Vr, (others=>'Z') after 1 ps;
XbG_V145<=(others=>'Z');
XbG_V146<=Vr, (others=>'Z') after 1 ps;
XbG_V147<=(others=>'Z');
XbG_V148<=Vr, (others=>'Z') after 1 ps;
XbG_V149<=(others=>'Z');
XbG_V15<=(others=>'Z');
XbG_V150<=Vr, (others=>'Z') after 1 ps;
XbG_V151<=(others=>'Z');
XbG_V152<=Vr, (others=>'Z') after 1 ps;
XbG_V153<=(others=>'Z');
XbG_V154<=Vr, (others=>'Z') after 1 ps;
XbG_V155<=(others=>'Z');
XbG_V156<=Vr, (others=>'Z') after 1 ps;
XbG_V157<=(others=>'Z');
XbG_V158<=Vr, (others=>'Z') after 1 ps;
XbG_V159<=(others=>'Z');
XbG_V16<=(others=>'Z');
XbG_V160<=Vr, (others=>'Z') after 1 ps;
XbG_V161<=(others=>'Z');
XbG_V162<=Vr, (others=>'Z') after 1 ps;
XbG_V163<=(others=>'Z');
XbG_V164<=Vr, (others=>'Z') after 1 ps;
XbG_V165<=(others=>'Z');
XbG_V166<=Vr, (others=>'Z') after 1 ps;
XbG_V167<=(others=>'Z');
XbG_V168<=Vr, (others=>'Z') after 1 ps;
XbG_V169<=(others=>'Z');
XbG_V17<=(others=>'Z');
XbG_V170<=Vr, (others=>'Z') after 1 ps;
XbG_V171<=(others=>'Z');
XbG_V172<=Vr, (others=>'Z') after 1 ps;
XbG_V173<=(others=>'Z');
XbG_V174<=Vr, (others=>'Z') after 1 ps;
XbG_V175<=(others=>'Z');
XbG_V176<=Vr, (others=>'Z') after 1 ps;
XbG_V177<=(others=>'Z');
XbG_V178<=Vr, (others=>'Z') after 1 ps;
XbG_V179<=(others=>'Z');
XbG_V18<=(others=>'Z');
XbG_V180<=Vr, (others=>'Z') after 1 ps;
XbG_V181<=(others=>'Z');
XbG_V182<=Vr, (others=>'Z') after 1 ps;
XbG_V183<=(others=>'Z');
XbG_V184<=Vr, (others=>'Z') after 1 ps;
XbG_V185<=(others=>'Z');
XbG_V186<=Vr, (others=>'Z') after 1 ps;
XbG_V187<=(others=>'Z');
XbG_V188<=Vr, (others=>'Z') after 1 ps;
XbG_V189<=(others=>'Z');
XbG_V19<=(others=>'Z');
XbG_V2<=(others=>'Z');
XbG_V20<=(others=>'Z');
XbG_V21<=(others=>'Z');
XbG_V22<=(others=>'Z');
XbG_V23<=(others=>'Z');
XbG_V24<=(others=>'Z');
XbG_V25<=(others=>'Z');
XbG_V26<=(others=>'Z');
XbG_V27<=(others=>'Z');
XbG_V28<=(others=>'Z');
XbG_V29<=(others=>'Z');
XbG_V3<=(others=>'Z');
XbG_V30<=(others=>'Z');
XbG_V31<=(others=>'Z');
XbG_V32<=(others=>'Z');
XbG_V33<=(others=>'Z');
XbG_V34<=(others=>'Z');
XbG_V35<=(others=>'Z');
XbG_V36<=(others=>'Z');
XbG_V37<=(others=>'Z');
XbG_V38<=(others=>'Z');
XbG_V39<=(others=>'Z');
XbG_V4<=(others=>'Z');
XbG_V40<=(others=>'Z');
XbG_V41<=(others=>'Z');
XbG_V42<=(others=>'Z');
XbG_V43<=(others=>'Z');
XbG_V44<=(others=>'Z');
XbG_V45<=(others=>'Z');
XbG_V46<=(others=>'Z');
XbG_V47<=(others=>'Z');
XbG_V48<=(others=>'Z');
XbG_V49<=(others=>'Z');
XbG_V5<=(others=>'Z');
XbG_V50<=(others=>'Z');
XbG_V51<=(others=>'Z');
XbG_V52<=(others=>'Z');
XbG_V53<=(others=>'Z');
XbG_V54<=(others=>'Z');
XbG_V55<=(others=>'Z');
XbG_V56<=(others=>'Z');
XbG_V57<=(others=>'Z');
XbG_V58<=(others=>'Z');
XbG_V59<=(others=>'Z');
XbG_V6<=(others=>'Z');
XbG_V60<=(others=>'Z');
XbG_V61<=(others=>'Z');
XbG_V62<=(others=>'Z');
XbG_V63<=(others=>'Z');
XbG_V64<=(others=>'Z');
XbG_V65<=(others=>'Z');
XbG_V66<=(others=>'Z');
XbG_V67<=(others=>'Z');
XbG_V68<=Vr, (others=>'Z') after 1 ps;
XbG_V69<=(others=>'Z');
XbG_V7<=(others=>'Z');
XbG_V70<=Vr, (others=>'Z') after 1 ps;
XbG_V71<=(others=>'Z');
XbG_V72<=Vr, (others=>'Z') after 1 ps;
XbG_V73<=(others=>'Z');
XbG_V74<=Vr, (others=>'Z') after 1 ps;
XbG_V75<=(others=>'Z');
XbG_V76<=Vr, (others=>'Z') after 1 ps;
XbG_V77<=(others=>'Z');
XbG_V78<=Vr, (others=>'Z') after 1 ps;
XbG_V79<=(others=>'Z');
XbG_V8<=(others=>'Z');
XbG_V80<=Vr, (others=>'Z') after 1 ps;
XbG_V81<=(others=>'Z');
XbG_V82<=Vr, (others=>'Z') after 1 ps;
XbG_V83<=(others=>'Z');
XbG_V84<=Vr, (others=>'Z') after 1 ps;
XbG_V85<=(others=>'Z');
XbG_V86<=Vr, (others=>'Z') after 1 ps;
XbG_V87<=(others=>'Z');
XbG_V88<=Vr, (others=>'Z') after 1 ps;
XbG_V89<=(others=>'Z');
XbG_V9<=(others=>'Z');
XbG_V90<=Vr, (others=>'Z') after 1 ps;
XbG_V91<=(others=>'Z');
XbG_V92<=Vr, (others=>'Z') after 1 ps;
XbG_V93<=(others=>'Z');
XbG_V94<=Vr, (others=>'Z') after 1 ps;
XbG_V95<=(others=>'Z');
XbG_V96<=Vr, (others=>'Z') after 1 ps;
XbG_V97<=(others=>'Z');
XbG_V98<=Vr, (others=>'Z') after 1 ps;
XbG_V99<=(others=>'Z');

done<='1' after clk_period;

feedback_enable <= '1';

next_state<=IDLE;

end case;

end process;

end Behavioral;
